library gp;
context gp.std_context;

package programs_tuples_nicolau_c_pkg is 

  constant opcode_type : type_t := uint_type(8);
  constant opcode_width : positive := get_width(opcode_type);

  constant programs : tuple_array(0 to 30)(0 to 4095)(7 downto 0) := (
    -- Bin `1`...
    0 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#B9#),
      1 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#0D#),
      33 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#0C#),
      65 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#0E#),
      97 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#0F#),
      129 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#0B#),
      161 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#11#),
      193 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#0A#),
      225 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#BF#),
      257 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#C4#),
      289 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#10#),
      321 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#2D#),
      353 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#4A#),
      385 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#8B#),
      417 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#C1#),
      449 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#92#),
      481 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#8A#),
      513 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#1F#),
      545 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#D3#),
      577 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#D4#),
      609 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#2F#),
      641 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#F2#),
      673 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#5F#),
      705 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#A5#),
      737 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#1D#),
      769 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#71#),
      801 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#B8#),
      833 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#30#),
      865 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#5B#),
      897 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#76#),
      929 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#61#),
      961 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#81#),
      993 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#CC#),
      1025 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#F4#),
      1057 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#9F#),
      1089 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#97#),
      1121 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#BB#),
      1153 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#85#),
      1185 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#7C#),
      1217 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#A2#),
      1249 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#69#),
      1281 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#46#),
      1313 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#DB#),
      1345 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#B0#),
      1377 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#B4#),
      1409 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#36#),
      1441 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#CE#),
      1473 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#9B#),
      1505 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#E7#),
      1537 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#B3#),
      1569 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#5D#),
      1601 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#D1#),
      1633 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#41#),
      1665 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#34#),
      1697 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#C5#),
      1729 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#64#),
      1761 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#B6#),
      1793 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#23#),
      1825 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#F1#),
      1857 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#98#),
      1889 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#E0#),
      1921 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#ED#),
      1953 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#E1#),
      1985 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#2C#),
      2017 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#9D#),
      2049 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#4E#),
      2081 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#59#),
      2113 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#DD#),
      2145 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#1A#),
      2177 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#82#),
      2209 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#2A#),
      2241 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#8F#),
      2273 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#26#),
      2305 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#FC#),
      2337 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#B7#),
      2369 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#91#),
      2401 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#DA#),
      2433 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#7A#),
      2465 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#1E#),
      2497 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#C3#),
      2529 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#AC#),
      2561 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#B2#),
      2593 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#29#),
      2625 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#BA#),
      2657 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#F7#),
      2689 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#EF#),
      2721 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#87#),
      2753 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#44#),
      2785 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#FB#),
      2817 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#60#),
      2849 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#72#),
      2881 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#49#),
      2913 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#4B#),
      2945 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#E8#),
      2977 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#AE#),
      3009 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#58#),
      3041 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#D6#),
      3073 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#9E#),
      3105 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#DF#),
      3137 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#39#),
      3169 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#6E#),
      3201 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#3D#),
      3233 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#D0#),
      3265 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#F6#),
      3297 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#18#),
      3329 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#80#),
      3361 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#32#),
      3393 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#9A#),
      3425 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#BD#),
      3457 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#DE#),
      3489 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#47#),
      3521 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#6D#),
      3553 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#AA#),
      3585 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#27#),
      3617 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#17#),
      3649 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#84#),
      3681 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#54#),
      3713 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#A0#),
      3745 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#96#),
      3777 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#68#),
      3809 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#D9#),
      3841 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#E4#),
      3873 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#8E#),
      3905 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#56#),
      3937 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#89#),
      3969 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#5E#),
      4001 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#C7#),
      4033 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#33#),
      4065 to 4095 => (others => '0')
  ),

    -- Bin `2`...
    1 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#01#),
      1 => to_slv(opcode_type, 16#0F#),
      2 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#01#),
      33 => to_slv(opcode_type, 16#9F#),
      34 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#04#),
      65 => to_slv(opcode_type, 16#0D#),
      66 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#02#),
      97 => to_slv(opcode_type, 16#0B#),
      98 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#05#),
      129 => to_slv(opcode_type, 16#0B#),
      130 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#03#),
      161 => to_slv(opcode_type, 16#0C#),
      162 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#03#),
      193 => to_slv(opcode_type, 16#0A#),
      194 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#04#),
      225 => to_slv(opcode_type, 16#0B#),
      226 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#02#),
      257 => to_slv(opcode_type, 16#51#),
      258 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#05#),
      289 => to_slv(opcode_type, 16#0F#),
      290 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#02#),
      321 => to_slv(opcode_type, 16#0E#),
      322 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#05#),
      353 => to_slv(opcode_type, 16#0E#),
      354 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#02#),
      385 => to_slv(opcode_type, 16#11#),
      386 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#01#),
      417 => to_slv(opcode_type, 16#10#),
      418 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#01#),
      449 => to_slv(opcode_type, 16#0E#),
      450 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#04#),
      481 => to_slv(opcode_type, 16#0C#),
      482 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#03#),
      513 => to_slv(opcode_type, 16#0D#),
      514 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#04#),
      545 => to_slv(opcode_type, 16#0F#),
      546 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#04#),
      577 => to_slv(opcode_type, 16#B5#),
      578 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#02#),
      609 => to_slv(opcode_type, 16#10#),
      610 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#05#),
      641 => to_slv(opcode_type, 16#0C#),
      642 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#02#),
      673 => to_slv(opcode_type, 16#0F#),
      674 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#04#),
      705 => to_slv(opcode_type, 16#58#),
      706 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#04#),
      737 => to_slv(opcode_type, 16#11#),
      738 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#04#),
      769 => to_slv(opcode_type, 16#0E#),
      770 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#03#),
      801 => to_slv(opcode_type, 16#0E#),
      802 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#02#),
      833 => to_slv(opcode_type, 16#73#),
      834 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#01#),
      865 => to_slv(opcode_type, 16#0C#),
      866 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#03#),
      897 => to_slv(opcode_type, 16#10#),
      898 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#02#),
      929 => to_slv(opcode_type, 16#0C#),
      930 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#05#),
      961 => to_slv(opcode_type, 16#0A#),
      962 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#01#),
      993 => to_slv(opcode_type, 16#0A#),
      994 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#05#),
      1025 => to_slv(opcode_type, 16#11#),
      1026 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#01#),
      1057 => to_slv(opcode_type, 16#0D#),
      1058 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#01#),
      1089 => to_slv(opcode_type, 16#11#),
      1090 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#04#),
      1121 => to_slv(opcode_type, 16#0A#),
      1122 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#01#),
      1153 => to_slv(opcode_type, 16#A1#),
      1154 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#02#),
      1185 => to_slv(opcode_type, 16#64#),
      1186 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#02#),
      1217 => to_slv(opcode_type, 16#0A#),
      1218 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#01#),
      1249 => to_slv(opcode_type, 16#0B#),
      1250 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#04#),
      1281 => to_slv(opcode_type, 16#10#),
      1282 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#02#),
      1313 => to_slv(opcode_type, 16#7F#),
      1314 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#05#),
      1345 => to_slv(opcode_type, 16#E3#),
      1346 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#05#),
      1377 => to_slv(opcode_type, 16#10#),
      1378 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#03#),
      1409 => to_slv(opcode_type, 16#43#),
      1410 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#03#),
      1441 => to_slv(opcode_type, 16#11#),
      1442 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#03#),
      1473 => to_slv(opcode_type, 16#0B#),
      1474 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#01#),
      1505 => to_slv(opcode_type, 16#70#),
      1506 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#03#),
      1537 => to_slv(opcode_type, 16#38#),
      1538 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#02#),
      1569 => to_slv(opcode_type, 16#D0#),
      1570 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#03#),
      1601 => to_slv(opcode_type, 16#52#),
      1602 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#05#),
      1633 => to_slv(opcode_type, 16#0D#),
      1634 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#03#),
      1665 => to_slv(opcode_type, 16#15#),
      1666 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#04#),
      1697 => to_slv(opcode_type, 16#8B#),
      1698 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#02#),
      1729 => to_slv(opcode_type, 16#0D#),
      1730 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#02#),
      1761 => to_slv(opcode_type, 16#FD#),
      1762 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#03#),
      1793 => to_slv(opcode_type, 16#FA#),
      1794 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#01#),
      1825 => to_slv(opcode_type, 16#53#),
      1826 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#04#),
      1857 => to_slv(opcode_type, 16#67#),
      1858 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#05#),
      1889 => to_slv(opcode_type, 16#50#),
      1890 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#05#),
      1921 => to_slv(opcode_type, 16#33#),
      1922 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#03#),
      1953 => to_slv(opcode_type, 16#0F#),
      1954 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#03#),
      1985 => to_slv(opcode_type, 16#F5#),
      1986 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#05#),
      2017 => to_slv(opcode_type, 16#B6#),
      2018 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#04#),
      2049 => to_slv(opcode_type, 16#86#),
      2050 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#04#),
      2081 => to_slv(opcode_type, 16#17#),
      2082 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#05#),
      2113 => to_slv(opcode_type, 16#59#),
      2114 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#01#),
      2145 => to_slv(opcode_type, 16#93#),
      2146 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#04#),
      2177 => to_slv(opcode_type, 16#8E#),
      2178 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#05#),
      2209 => to_slv(opcode_type, 16#3D#),
      2210 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#01#),
      2241 => to_slv(opcode_type, 16#FC#),
      2242 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#03#),
      2273 => to_slv(opcode_type, 16#41#),
      2274 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#05#),
      2305 => to_slv(opcode_type, 16#A6#),
      2306 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#01#),
      2337 => to_slv(opcode_type, 16#B5#),
      2338 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#04#),
      2369 => to_slv(opcode_type, 16#D8#),
      2370 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#04#),
      2401 => to_slv(opcode_type, 16#6A#),
      2402 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#05#),
      2433 => to_slv(opcode_type, 16#43#),
      2434 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#03#),
      2465 => to_slv(opcode_type, 16#49#),
      2466 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#01#),
      2497 => to_slv(opcode_type, 16#4C#),
      2498 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#02#),
      2529 => to_slv(opcode_type, 16#5D#),
      2530 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#01#),
      2561 => to_slv(opcode_type, 16#CD#),
      2562 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#01#),
      2593 => to_slv(opcode_type, 16#3E#),
      2594 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#04#),
      2625 => to_slv(opcode_type, 16#49#),
      2626 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#04#),
      2657 => to_slv(opcode_type, 16#64#),
      2658 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#02#),
      2689 => to_slv(opcode_type, 16#1F#),
      2690 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#02#),
      2721 => to_slv(opcode_type, 16#7A#),
      2722 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#02#),
      2753 => to_slv(opcode_type, 16#CE#),
      2754 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#01#),
      2785 => to_slv(opcode_type, 16#51#),
      2786 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#01#),
      2817 => to_slv(opcode_type, 16#22#),
      2818 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#02#),
      2849 => to_slv(opcode_type, 16#9E#),
      2850 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#05#),
      2881 => to_slv(opcode_type, 16#42#),
      2882 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#01#),
      2913 => to_slv(opcode_type, 16#E3#),
      2914 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#04#),
      2945 => to_slv(opcode_type, 16#1E#),
      2946 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#03#),
      2977 => to_slv(opcode_type, 16#2B#),
      2978 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#04#),
      3009 => to_slv(opcode_type, 16#46#),
      3010 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#02#),
      3041 => to_slv(opcode_type, 16#5B#),
      3042 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#05#),
      3073 => to_slv(opcode_type, 16#5E#),
      3074 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#03#),
      3105 => to_slv(opcode_type, 16#7B#),
      3106 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#04#),
      3137 => to_slv(opcode_type, 16#1A#),
      3138 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#02#),
      3169 => to_slv(opcode_type, 16#EC#),
      3170 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#03#),
      3201 => to_slv(opcode_type, 16#A5#),
      3202 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#01#),
      3233 => to_slv(opcode_type, 16#EB#),
      3234 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#02#),
      3265 => to_slv(opcode_type, 16#43#),
      3266 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#01#),
      3297 => to_slv(opcode_type, 16#9C#),
      3298 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#01#),
      3329 => to_slv(opcode_type, 16#66#),
      3330 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#01#),
      3361 => to_slv(opcode_type, 16#D0#),
      3362 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#05#),
      3393 => to_slv(opcode_type, 16#9E#),
      3394 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#04#),
      3425 => to_slv(opcode_type, 16#39#),
      3426 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#02#),
      3457 => to_slv(opcode_type, 16#3C#),
      3458 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#03#),
      3489 => to_slv(opcode_type, 16#92#),
      3490 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#02#),
      3521 => to_slv(opcode_type, 16#52#),
      3522 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#02#),
      3553 => to_slv(opcode_type, 16#96#),
      3554 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#01#),
      3585 => to_slv(opcode_type, 16#F5#),
      3586 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#05#),
      3617 => to_slv(opcode_type, 16#B0#),
      3618 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#05#),
      3649 => to_slv(opcode_type, 16#D0#),
      3650 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#04#),
      3681 => to_slv(opcode_type, 16#1C#),
      3682 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#04#),
      3713 => to_slv(opcode_type, 16#AA#),
      3714 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#02#),
      3745 => to_slv(opcode_type, 16#1B#),
      3746 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#05#),
      3777 => to_slv(opcode_type, 16#56#),
      3778 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#05#),
      3809 => to_slv(opcode_type, 16#CA#),
      3810 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#01#),
      3841 => to_slv(opcode_type, 16#EF#),
      3842 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#04#),
      3873 => to_slv(opcode_type, 16#18#),
      3874 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#03#),
      3905 => to_slv(opcode_type, 16#35#),
      3906 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#03#),
      3937 => to_slv(opcode_type, 16#95#),
      3938 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#04#),
      3969 => to_slv(opcode_type, 16#84#),
      3970 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#01#),
      4001 => to_slv(opcode_type, 16#AA#),
      4002 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#02#),
      4033 => to_slv(opcode_type, 16#CB#),
      4034 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#05#),
      4065 => to_slv(opcode_type, 16#B8#),
      4066 to 4095 => (others => '0')
  ),

    -- Bin `3`...
    2 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#09#),
      1 => to_slv(opcode_type, 16#0D#),
      2 => to_slv(opcode_type, 16#0E#),
      3 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#02#),
      33 => to_slv(opcode_type, 16#01#),
      34 => to_slv(opcode_type, 16#0B#),
      35 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#07#),
      65 => to_slv(opcode_type, 16#10#),
      66 => to_slv(opcode_type, 16#0D#),
      67 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#04#),
      97 => to_slv(opcode_type, 16#02#),
      98 => to_slv(opcode_type, 16#10#),
      99 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#04#),
      129 => to_slv(opcode_type, 16#01#),
      130 => to_slv(opcode_type, 16#0B#),
      131 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#03#),
      161 => to_slv(opcode_type, 16#01#),
      162 => to_slv(opcode_type, 16#0D#),
      163 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#06#),
      193 => to_slv(opcode_type, 16#10#),
      194 => to_slv(opcode_type, 16#0A#),
      195 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#03#),
      225 => to_slv(opcode_type, 16#03#),
      226 => to_slv(opcode_type, 16#10#),
      227 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#07#),
      257 => to_slv(opcode_type, 16#0D#),
      258 => to_slv(opcode_type, 16#0A#),
      259 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#51#),
      290 => to_slv(opcode_type, 16#0E#),
      291 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#02#),
      321 => to_slv(opcode_type, 16#02#),
      322 => to_slv(opcode_type, 16#0A#),
      323 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#03#),
      353 => to_slv(opcode_type, 16#03#),
      354 => to_slv(opcode_type, 16#0B#),
      355 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#04#),
      385 => to_slv(opcode_type, 16#05#),
      386 => to_slv(opcode_type, 16#10#),
      387 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#09#),
      417 => to_slv(opcode_type, 16#0E#),
      418 => to_slv(opcode_type, 16#0D#),
      419 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#06#),
      449 => to_slv(opcode_type, 16#0A#),
      450 => to_slv(opcode_type, 16#0F#),
      451 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#01#),
      481 => to_slv(opcode_type, 16#05#),
      482 => to_slv(opcode_type, 16#0C#),
      483 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#03#),
      513 => to_slv(opcode_type, 16#05#),
      514 => to_slv(opcode_type, 16#11#),
      515 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#02#),
      545 => to_slv(opcode_type, 16#02#),
      546 => to_slv(opcode_type, 16#11#),
      547 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#01#),
      577 => to_slv(opcode_type, 16#05#),
      578 => to_slv(opcode_type, 16#94#),
      579 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#06#),
      609 => to_slv(opcode_type, 16#0D#),
      610 => to_slv(opcode_type, 16#0D#),
      611 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#02#),
      641 => to_slv(opcode_type, 16#01#),
      642 => to_slv(opcode_type, 16#FF#),
      643 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#06#),
      673 => to_slv(opcode_type, 16#0A#),
      674 => to_slv(opcode_type, 16#11#),
      675 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#06#),
      705 => to_slv(opcode_type, 16#10#),
      706 => to_slv(opcode_type, 16#0F#),
      707 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#09#),
      737 => to_slv(opcode_type, 16#0F#),
      738 => to_slv(opcode_type, 16#0A#),
      739 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#01#),
      769 => to_slv(opcode_type, 16#01#),
      770 => to_slv(opcode_type, 16#10#),
      771 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#06#),
      801 => to_slv(opcode_type, 16#0E#),
      802 => to_slv(opcode_type, 16#10#),
      803 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#02#),
      833 => to_slv(opcode_type, 16#05#),
      834 => to_slv(opcode_type, 16#0E#),
      835 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#04#),
      865 => to_slv(opcode_type, 16#04#),
      866 => to_slv(opcode_type, 16#A8#),
      867 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#08#),
      897 => to_slv(opcode_type, 16#0B#),
      898 => to_slv(opcode_type, 16#11#),
      899 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#04#),
      929 => to_slv(opcode_type, 16#04#),
      930 => to_slv(opcode_type, 16#0F#),
      931 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#11#),
      962 => to_slv(opcode_type, 16#0E#),
      963 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#09#),
      993 => to_slv(opcode_type, 16#10#),
      994 => to_slv(opcode_type, 16#D9#),
      995 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#05#),
      1025 => to_slv(opcode_type, 16#05#),
      1026 => to_slv(opcode_type, 16#10#),
      1027 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#03#),
      1057 => to_slv(opcode_type, 16#04#),
      1058 => to_slv(opcode_type, 16#0B#),
      1059 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#09#),
      1089 => to_slv(opcode_type, 16#0E#),
      1090 => to_slv(opcode_type, 16#11#),
      1091 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#01#),
      1121 => to_slv(opcode_type, 16#03#),
      1122 => to_slv(opcode_type, 16#0E#),
      1123 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#01#),
      1153 => to_slv(opcode_type, 16#03#),
      1154 => to_slv(opcode_type, 16#0F#),
      1155 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#03#),
      1185 => to_slv(opcode_type, 16#02#),
      1186 => to_slv(opcode_type, 16#0A#),
      1187 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#05#),
      1217 => to_slv(opcode_type, 16#02#),
      1218 => to_slv(opcode_type, 16#0F#),
      1219 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#03#),
      1249 => to_slv(opcode_type, 16#03#),
      1250 => to_slv(opcode_type, 16#0C#),
      1251 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#0C#),
      1282 => to_slv(opcode_type, 16#0F#),
      1283 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#02#),
      1313 => to_slv(opcode_type, 16#05#),
      1314 => to_slv(opcode_type, 16#EB#),
      1315 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#04#),
      1345 => to_slv(opcode_type, 16#04#),
      1346 => to_slv(opcode_type, 16#0B#),
      1347 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#03#),
      1377 => to_slv(opcode_type, 16#05#),
      1378 => to_slv(opcode_type, 16#0E#),
      1379 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#F5#),
      1410 => to_slv(opcode_type, 16#0E#),
      1411 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#05#),
      1441 => to_slv(opcode_type, 16#02#),
      1442 => to_slv(opcode_type, 16#10#),
      1443 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#04#),
      1473 => to_slv(opcode_type, 16#02#),
      1474 => to_slv(opcode_type, 16#0D#),
      1475 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#02#),
      1505 => to_slv(opcode_type, 16#03#),
      1506 => to_slv(opcode_type, 16#0B#),
      1507 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#09#),
      1537 => to_slv(opcode_type, 16#0E#),
      1538 => to_slv(opcode_type, 16#0A#),
      1539 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#03#),
      1569 => to_slv(opcode_type, 16#05#),
      1570 => to_slv(opcode_type, 16#0D#),
      1571 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#02#),
      1601 => to_slv(opcode_type, 16#05#),
      1602 => to_slv(opcode_type, 16#0C#),
      1603 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#01#),
      1633 => to_slv(opcode_type, 16#03#),
      1634 => to_slv(opcode_type, 16#0A#),
      1635 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#0C#),
      1666 => to_slv(opcode_type, 16#0E#),
      1667 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#06#),
      1697 => to_slv(opcode_type, 16#10#),
      1698 => to_slv(opcode_type, 16#11#),
      1699 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#04#),
      1729 => to_slv(opcode_type, 16#02#),
      1730 => to_slv(opcode_type, 16#0F#),
      1731 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#03#),
      1761 => to_slv(opcode_type, 16#04#),
      1762 => to_slv(opcode_type, 16#0A#),
      1763 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#04#),
      1793 => to_slv(opcode_type, 16#05#),
      1794 => to_slv(opcode_type, 16#BD#),
      1795 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#01#),
      1825 => to_slv(opcode_type, 16#02#),
      1826 => to_slv(opcode_type, 16#0B#),
      1827 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#08#),
      1857 => to_slv(opcode_type, 16#11#),
      1858 => to_slv(opcode_type, 16#0A#),
      1859 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#04#),
      1889 => to_slv(opcode_type, 16#04#),
      1890 => to_slv(opcode_type, 16#11#),
      1891 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#07#),
      1921 => to_slv(opcode_type, 16#0E#),
      1922 => to_slv(opcode_type, 16#0A#),
      1923 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#08#),
      1953 => to_slv(opcode_type, 16#0F#),
      1954 => to_slv(opcode_type, 16#0B#),
      1955 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#02#),
      1985 => to_slv(opcode_type, 16#02#),
      1986 => to_slv(opcode_type, 16#10#),
      1987 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#09#),
      2017 => to_slv(opcode_type, 16#0C#),
      2018 => to_slv(opcode_type, 16#10#),
      2019 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#01#),
      2049 => to_slv(opcode_type, 16#01#),
      2050 => to_slv(opcode_type, 16#0E#),
      2051 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#07#),
      2081 => to_slv(opcode_type, 16#0F#),
      2082 => to_slv(opcode_type, 16#0E#),
      2083 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#02#),
      2113 => to_slv(opcode_type, 16#05#),
      2114 => to_slv(opcode_type, 16#0B#),
      2115 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#01#),
      2145 => to_slv(opcode_type, 16#02#),
      2146 => to_slv(opcode_type, 16#0E#),
      2147 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#03#),
      2177 => to_slv(opcode_type, 16#04#),
      2178 => to_slv(opcode_type, 16#11#),
      2179 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#01#),
      2209 => to_slv(opcode_type, 16#02#),
      2210 => to_slv(opcode_type, 16#11#),
      2211 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#0D#),
      2242 => to_slv(opcode_type, 16#A8#),
      2243 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#02#),
      2273 => to_slv(opcode_type, 16#04#),
      2274 => to_slv(opcode_type, 16#10#),
      2275 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#08#),
      2305 => to_slv(opcode_type, 16#0F#),
      2306 => to_slv(opcode_type, 16#0E#),
      2307 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#03#),
      2337 => to_slv(opcode_type, 16#05#),
      2338 => to_slv(opcode_type, 16#0F#),
      2339 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#09#),
      2369 => to_slv(opcode_type, 16#0E#),
      2370 => to_slv(opcode_type, 16#0C#),
      2371 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#09#),
      2401 => to_slv(opcode_type, 16#0D#),
      2402 => to_slv(opcode_type, 16#0C#),
      2403 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#07#),
      2433 => to_slv(opcode_type, 16#0E#),
      2434 => to_slv(opcode_type, 16#0C#),
      2435 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#02#),
      2465 => to_slv(opcode_type, 16#01#),
      2466 => to_slv(opcode_type, 16#0D#),
      2467 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#05#),
      2497 => to_slv(opcode_type, 16#04#),
      2498 => to_slv(opcode_type, 16#0A#),
      2499 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#F2#),
      2530 => to_slv(opcode_type, 16#0E#),
      2531 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#01#),
      2561 => to_slv(opcode_type, 16#05#),
      2562 => to_slv(opcode_type, 16#0F#),
      2563 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#05#),
      2593 => to_slv(opcode_type, 16#05#),
      2594 => to_slv(opcode_type, 16#11#),
      2595 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#08#),
      2625 => to_slv(opcode_type, 16#11#),
      2626 => to_slv(opcode_type, 16#0F#),
      2627 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#06#),
      2657 => to_slv(opcode_type, 16#11#),
      2658 => to_slv(opcode_type, 16#0B#),
      2659 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#02#),
      2689 => to_slv(opcode_type, 16#01#),
      2690 => to_slv(opcode_type, 16#3C#),
      2691 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#03#),
      2721 => to_slv(opcode_type, 16#01#),
      2722 => to_slv(opcode_type, 16#0E#),
      2723 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#09#),
      2753 => to_slv(opcode_type, 16#11#),
      2754 => to_slv(opcode_type, 16#DA#),
      2755 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#02#),
      2785 => to_slv(opcode_type, 16#05#),
      2786 => to_slv(opcode_type, 16#10#),
      2787 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#02#),
      2817 => to_slv(opcode_type, 16#03#),
      2818 => to_slv(opcode_type, 16#0A#),
      2819 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#08#),
      2849 => to_slv(opcode_type, 16#10#),
      2850 => to_slv(opcode_type, 16#0D#),
      2851 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#02#),
      2881 => to_slv(opcode_type, 16#05#),
      2882 => to_slv(opcode_type, 16#0F#),
      2883 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#01#),
      2913 => to_slv(opcode_type, 16#04#),
      2914 => to_slv(opcode_type, 16#0D#),
      2915 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#08#),
      2945 => to_slv(opcode_type, 16#0C#),
      2946 => to_slv(opcode_type, 16#0B#),
      2947 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#07#),
      2977 => to_slv(opcode_type, 16#0B#),
      2978 => to_slv(opcode_type, 16#0C#),
      2979 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#01#),
      3009 => to_slv(opcode_type, 16#01#),
      3010 => to_slv(opcode_type, 16#84#),
      3011 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#06#),
      3041 => to_slv(opcode_type, 16#11#),
      3042 => to_slv(opcode_type, 16#10#),
      3043 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#05#),
      3073 => to_slv(opcode_type, 16#03#),
      3074 => to_slv(opcode_type, 16#0D#),
      3075 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#06#),
      3105 => to_slv(opcode_type, 16#0B#),
      3106 => to_slv(opcode_type, 16#0A#),
      3107 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#09#),
      3137 => to_slv(opcode_type, 16#0E#),
      3138 => to_slv(opcode_type, 16#0F#),
      3139 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#04#),
      3169 => to_slv(opcode_type, 16#04#),
      3170 => to_slv(opcode_type, 16#0A#),
      3171 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#05#),
      3201 => to_slv(opcode_type, 16#04#),
      3202 => to_slv(opcode_type, 16#AF#),
      3203 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#0A#),
      3234 => to_slv(opcode_type, 16#0D#),
      3235 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#07#),
      3265 => to_slv(opcode_type, 16#0C#),
      3266 => to_slv(opcode_type, 16#0C#),
      3267 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#05#),
      3297 => to_slv(opcode_type, 16#05#),
      3298 => to_slv(opcode_type, 16#0B#),
      3299 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#04#),
      3329 => to_slv(opcode_type, 16#04#),
      3330 => to_slv(opcode_type, 16#10#),
      3331 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#06#),
      3361 => to_slv(opcode_type, 16#0B#),
      3362 => to_slv(opcode_type, 16#0D#),
      3363 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#08#),
      3393 => to_slv(opcode_type, 16#11#),
      3394 => to_slv(opcode_type, 16#10#),
      3395 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#01#),
      3425 => to_slv(opcode_type, 16#04#),
      3426 => to_slv(opcode_type, 16#0E#),
      3427 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#07#),
      3457 => to_slv(opcode_type, 16#0D#),
      3458 => to_slv(opcode_type, 16#11#),
      3459 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#06#),
      3489 => to_slv(opcode_type, 16#0A#),
      3490 => to_slv(opcode_type, 16#7A#),
      3491 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#09#),
      3521 => to_slv(opcode_type, 16#0C#),
      3522 => to_slv(opcode_type, 16#0A#),
      3523 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#05#),
      3553 => to_slv(opcode_type, 16#02#),
      3554 => to_slv(opcode_type, 16#11#),
      3555 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#03#),
      3585 => to_slv(opcode_type, 16#05#),
      3586 => to_slv(opcode_type, 16#10#),
      3587 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#06#),
      3617 => to_slv(opcode_type, 16#0F#),
      3618 => to_slv(opcode_type, 16#0F#),
      3619 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#02#),
      3649 => to_slv(opcode_type, 16#02#),
      3650 => to_slv(opcode_type, 16#0C#),
      3651 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#05#),
      3681 => to_slv(opcode_type, 16#01#),
      3682 => to_slv(opcode_type, 16#0C#),
      3683 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#05#),
      3713 => to_slv(opcode_type, 16#01#),
      3714 => to_slv(opcode_type, 16#89#),
      3715 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#08#),
      3745 => to_slv(opcode_type, 16#0D#),
      3746 => to_slv(opcode_type, 16#2E#),
      3747 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#08#),
      3777 => to_slv(opcode_type, 16#0A#),
      3778 => to_slv(opcode_type, 16#70#),
      3779 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#02#),
      3809 => to_slv(opcode_type, 16#02#),
      3810 => to_slv(opcode_type, 16#0E#),
      3811 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#09#),
      3841 => to_slv(opcode_type, 16#0B#),
      3842 => to_slv(opcode_type, 16#0F#),
      3843 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#06#),
      3873 => to_slv(opcode_type, 16#0D#),
      3874 => to_slv(opcode_type, 16#11#),
      3875 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#02#),
      3905 => to_slv(opcode_type, 16#01#),
      3906 => to_slv(opcode_type, 16#0C#),
      3907 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#09#),
      3937 => to_slv(opcode_type, 16#10#),
      3938 => to_slv(opcode_type, 16#0C#),
      3939 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#01#),
      3969 => to_slv(opcode_type, 16#02#),
      3970 => to_slv(opcode_type, 16#10#),
      3971 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#08#),
      4001 => to_slv(opcode_type, 16#0C#),
      4002 => to_slv(opcode_type, 16#0C#),
      4003 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#04#),
      4033 => to_slv(opcode_type, 16#03#),
      4034 => to_slv(opcode_type, 16#0E#),
      4035 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#07#),
      4065 => to_slv(opcode_type, 16#21#),
      4066 => to_slv(opcode_type, 16#0E#),
      4067 to 4095 => (others => '0')
  ),

    -- Bin `4`...
    3 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#01#),
      1 => to_slv(opcode_type, 16#06#),
      2 => to_slv(opcode_type, 16#9C#),
      3 => to_slv(opcode_type, 16#13#),
      4 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#03#),
      33 => to_slv(opcode_type, 16#05#),
      34 => to_slv(opcode_type, 16#01#),
      35 => to_slv(opcode_type, 16#3A#),
      36 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#03#),
      65 => to_slv(opcode_type, 16#09#),
      66 => to_slv(opcode_type, 16#0B#),
      67 => to_slv(opcode_type, 16#0E#),
      68 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#07#),
      97 => to_slv(opcode_type, 16#03#),
      98 => to_slv(opcode_type, 16#0C#),
      99 => to_slv(opcode_type, 16#10#),
      100 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#01#),
      129 => to_slv(opcode_type, 16#01#),
      130 => to_slv(opcode_type, 16#05#),
      131 => to_slv(opcode_type, 16#0F#),
      132 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#01#),
      161 => to_slv(opcode_type, 16#05#),
      162 => to_slv(opcode_type, 16#05#),
      163 => to_slv(opcode_type, 16#0E#),
      164 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#05#),
      193 => to_slv(opcode_type, 16#02#),
      194 => to_slv(opcode_type, 16#02#),
      195 => to_slv(opcode_type, 16#62#),
      196 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#07#),
      225 => to_slv(opcode_type, 16#01#),
      226 => to_slv(opcode_type, 16#1D#),
      227 => to_slv(opcode_type, 16#0B#),
      228 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#09#),
      257 => to_slv(opcode_type, 16#05#),
      258 => to_slv(opcode_type, 16#0F#),
      259 => to_slv(opcode_type, 16#0F#),
      260 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#01#),
      289 => to_slv(opcode_type, 16#09#),
      290 => to_slv(opcode_type, 16#11#),
      291 => to_slv(opcode_type, 16#11#),
      292 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#03#),
      321 => to_slv(opcode_type, 16#04#),
      322 => to_slv(opcode_type, 16#02#),
      323 => to_slv(opcode_type, 16#10#),
      324 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#04#),
      353 => to_slv(opcode_type, 16#01#),
      354 => to_slv(opcode_type, 16#05#),
      355 => to_slv(opcode_type, 16#11#),
      356 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#08#),
      385 => to_slv(opcode_type, 16#03#),
      386 => to_slv(opcode_type, 16#0E#),
      387 => to_slv(opcode_type, 16#0F#),
      388 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#09#),
      417 => to_slv(opcode_type, 16#05#),
      418 => to_slv(opcode_type, 16#0D#),
      419 => to_slv(opcode_type, 16#0D#),
      420 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#06#),
      449 => to_slv(opcode_type, 16#01#),
      450 => to_slv(opcode_type, 16#0D#),
      451 => to_slv(opcode_type, 16#0E#),
      452 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#09#),
      481 => to_slv(opcode_type, 16#01#),
      482 => to_slv(opcode_type, 16#11#),
      483 => to_slv(opcode_type, 16#0E#),
      484 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#03#),
      514 => to_slv(opcode_type, 16#11#),
      515 => to_slv(opcode_type, 16#0A#),
      516 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#04#),
      545 => to_slv(opcode_type, 16#03#),
      546 => to_slv(opcode_type, 16#05#),
      547 => to_slv(opcode_type, 16#A7#),
      548 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#06#),
      577 => to_slv(opcode_type, 16#01#),
      578 => to_slv(opcode_type, 16#0B#),
      579 => to_slv(opcode_type, 16#9B#),
      580 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#06#),
      609 => to_slv(opcode_type, 16#03#),
      610 => to_slv(opcode_type, 16#0F#),
      611 => to_slv(opcode_type, 16#0E#),
      612 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#07#),
      641 => to_slv(opcode_type, 16#01#),
      642 => to_slv(opcode_type, 16#0C#),
      643 => to_slv(opcode_type, 16#0B#),
      644 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#01#),
      673 => to_slv(opcode_type, 16#09#),
      674 => to_slv(opcode_type, 16#10#),
      675 => to_slv(opcode_type, 16#26#),
      676 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#04#),
      705 => to_slv(opcode_type, 16#08#),
      706 => to_slv(opcode_type, 16#11#),
      707 => to_slv(opcode_type, 16#E7#),
      708 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#03#),
      737 => to_slv(opcode_type, 16#05#),
      738 => to_slv(opcode_type, 16#02#),
      739 => to_slv(opcode_type, 16#0C#),
      740 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#08#),
      769 => to_slv(opcode_type, 16#03#),
      770 => to_slv(opcode_type, 16#0A#),
      771 => to_slv(opcode_type, 16#0F#),
      772 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#08#),
      801 => to_slv(opcode_type, 16#03#),
      802 => to_slv(opcode_type, 16#0D#),
      803 => to_slv(opcode_type, 16#0E#),
      804 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#06#),
      833 => to_slv(opcode_type, 16#01#),
      834 => to_slv(opcode_type, 16#0F#),
      835 => to_slv(opcode_type, 16#0F#),
      836 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#01#),
      865 => to_slv(opcode_type, 16#03#),
      866 => to_slv(opcode_type, 16#03#),
      867 => to_slv(opcode_type, 16#0D#),
      868 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#08#),
      897 => to_slv(opcode_type, 16#03#),
      898 => to_slv(opcode_type, 16#0F#),
      899 => to_slv(opcode_type, 16#0E#),
      900 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#04#),
      929 => to_slv(opcode_type, 16#01#),
      930 => to_slv(opcode_type, 16#04#),
      931 => to_slv(opcode_type, 16#0E#),
      932 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#08#),
      961 => to_slv(opcode_type, 16#05#),
      962 => to_slv(opcode_type, 16#11#),
      963 => to_slv(opcode_type, 16#10#),
      964 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#03#),
      993 => to_slv(opcode_type, 16#01#),
      994 => to_slv(opcode_type, 16#05#),
      995 => to_slv(opcode_type, 16#0C#),
      996 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#09#),
      1025 => to_slv(opcode_type, 16#04#),
      1026 => to_slv(opcode_type, 16#10#),
      1027 => to_slv(opcode_type, 16#0C#),
      1028 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#08#),
      1057 => to_slv(opcode_type, 16#02#),
      1058 => to_slv(opcode_type, 16#0B#),
      1059 => to_slv(opcode_type, 16#0C#),
      1060 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#04#),
      1089 => to_slv(opcode_type, 16#07#),
      1090 => to_slv(opcode_type, 16#0F#),
      1091 => to_slv(opcode_type, 16#10#),
      1092 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#05#),
      1121 => to_slv(opcode_type, 16#04#),
      1122 => to_slv(opcode_type, 16#01#),
      1123 => to_slv(opcode_type, 16#10#),
      1124 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#05#),
      1153 => to_slv(opcode_type, 16#04#),
      1154 => to_slv(opcode_type, 16#02#),
      1155 => to_slv(opcode_type, 16#10#),
      1156 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#09#),
      1185 => to_slv(opcode_type, 16#05#),
      1186 => to_slv(opcode_type, 16#11#),
      1187 => to_slv(opcode_type, 16#0A#),
      1188 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#06#),
      1217 => to_slv(opcode_type, 16#05#),
      1218 => to_slv(opcode_type, 16#11#),
      1219 => to_slv(opcode_type, 16#0C#),
      1220 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#05#),
      1249 => to_slv(opcode_type, 16#07#),
      1250 => to_slv(opcode_type, 16#0B#),
      1251 => to_slv(opcode_type, 16#0F#),
      1252 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#07#),
      1281 => to_slv(opcode_type, 16#04#),
      1282 => to_slv(opcode_type, 16#10#),
      1283 => to_slv(opcode_type, 16#0F#),
      1284 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#02#),
      1313 => to_slv(opcode_type, 16#06#),
      1314 => to_slv(opcode_type, 16#10#),
      1315 => to_slv(opcode_type, 16#11#),
      1316 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#03#),
      1345 => to_slv(opcode_type, 16#03#),
      1346 => to_slv(opcode_type, 16#05#),
      1347 => to_slv(opcode_type, 16#C0#),
      1348 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#09#),
      1377 => to_slv(opcode_type, 16#01#),
      1378 => to_slv(opcode_type, 16#0D#),
      1379 => to_slv(opcode_type, 16#0A#),
      1380 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#01#),
      1409 => to_slv(opcode_type, 16#02#),
      1410 => to_slv(opcode_type, 16#01#),
      1411 => to_slv(opcode_type, 16#0A#),
      1412 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#08#),
      1441 => to_slv(opcode_type, 16#05#),
      1442 => to_slv(opcode_type, 16#11#),
      1443 => to_slv(opcode_type, 16#0F#),
      1444 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#03#),
      1473 => to_slv(opcode_type, 16#04#),
      1474 => to_slv(opcode_type, 16#05#),
      1475 => to_slv(opcode_type, 16#0E#),
      1476 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#06#),
      1505 => to_slv(opcode_type, 16#04#),
      1506 => to_slv(opcode_type, 16#0B#),
      1507 => to_slv(opcode_type, 16#0D#),
      1508 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#01#),
      1537 => to_slv(opcode_type, 16#01#),
      1538 => to_slv(opcode_type, 16#03#),
      1539 => to_slv(opcode_type, 16#0A#),
      1540 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#01#),
      1569 => to_slv(opcode_type, 16#03#),
      1570 => to_slv(opcode_type, 16#01#),
      1571 => to_slv(opcode_type, 16#9D#),
      1572 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#08#),
      1601 => to_slv(opcode_type, 16#04#),
      1602 => to_slv(opcode_type, 16#0F#),
      1603 => to_slv(opcode_type, 16#F0#),
      1604 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#06#),
      1633 => to_slv(opcode_type, 16#02#),
      1634 => to_slv(opcode_type, 16#10#),
      1635 => to_slv(opcode_type, 16#0E#),
      1636 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#07#),
      1665 => to_slv(opcode_type, 16#04#),
      1666 => to_slv(opcode_type, 16#10#),
      1667 => to_slv(opcode_type, 16#11#),
      1668 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#01#),
      1697 => to_slv(opcode_type, 16#05#),
      1698 => to_slv(opcode_type, 16#04#),
      1699 => to_slv(opcode_type, 16#0C#),
      1700 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#08#),
      1729 => to_slv(opcode_type, 16#05#),
      1730 => to_slv(opcode_type, 16#49#),
      1731 => to_slv(opcode_type, 16#10#),
      1732 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#06#),
      1761 => to_slv(opcode_type, 16#02#),
      1762 => to_slv(opcode_type, 16#0B#),
      1763 => to_slv(opcode_type, 16#0B#),
      1764 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#08#),
      1793 => to_slv(opcode_type, 16#05#),
      1794 => to_slv(opcode_type, 16#0A#),
      1795 => to_slv(opcode_type, 16#0C#),
      1796 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#02#),
      1825 => to_slv(opcode_type, 16#06#),
      1826 => to_slv(opcode_type, 16#0C#),
      1827 => to_slv(opcode_type, 16#10#),
      1828 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#01#),
      1857 => to_slv(opcode_type, 16#08#),
      1858 => to_slv(opcode_type, 16#9F#),
      1859 => to_slv(opcode_type, 16#0B#),
      1860 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#09#),
      1889 => to_slv(opcode_type, 16#04#),
      1890 => to_slv(opcode_type, 16#0E#),
      1891 => to_slv(opcode_type, 16#7C#),
      1892 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#05#),
      1921 => to_slv(opcode_type, 16#08#),
      1922 => to_slv(opcode_type, 16#8F#),
      1923 => to_slv(opcode_type, 16#BC#),
      1924 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#06#),
      1953 => to_slv(opcode_type, 16#02#),
      1954 => to_slv(opcode_type, 16#10#),
      1955 => to_slv(opcode_type, 16#0D#),
      1956 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#07#),
      1985 => to_slv(opcode_type, 16#04#),
      1986 => to_slv(opcode_type, 16#10#),
      1987 => to_slv(opcode_type, 16#10#),
      1988 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#01#),
      2017 => to_slv(opcode_type, 16#01#),
      2018 => to_slv(opcode_type, 16#03#),
      2019 => to_slv(opcode_type, 16#0F#),
      2020 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#02#),
      2049 => to_slv(opcode_type, 16#03#),
      2050 => to_slv(opcode_type, 16#02#),
      2051 => to_slv(opcode_type, 16#0A#),
      2052 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#07#),
      2081 => to_slv(opcode_type, 16#04#),
      2082 => to_slv(opcode_type, 16#0F#),
      2083 => to_slv(opcode_type, 16#0F#),
      2084 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#08#),
      2113 => to_slv(opcode_type, 16#03#),
      2114 => to_slv(opcode_type, 16#0E#),
      2115 => to_slv(opcode_type, 16#10#),
      2116 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#06#),
      2145 => to_slv(opcode_type, 16#03#),
      2146 => to_slv(opcode_type, 16#0F#),
      2147 => to_slv(opcode_type, 16#11#),
      2148 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#04#),
      2177 => to_slv(opcode_type, 16#05#),
      2178 => to_slv(opcode_type, 16#01#),
      2179 => to_slv(opcode_type, 16#0D#),
      2180 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#05#),
      2209 => to_slv(opcode_type, 16#08#),
      2210 => to_slv(opcode_type, 16#0D#),
      2211 => to_slv(opcode_type, 16#0E#),
      2212 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#07#),
      2241 => to_slv(opcode_type, 16#04#),
      2242 => to_slv(opcode_type, 16#0A#),
      2243 => to_slv(opcode_type, 16#0A#),
      2244 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#01#),
      2273 => to_slv(opcode_type, 16#01#),
      2274 => to_slv(opcode_type, 16#05#),
      2275 => to_slv(opcode_type, 16#0E#),
      2276 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#04#),
      2305 => to_slv(opcode_type, 16#07#),
      2306 => to_slv(opcode_type, 16#11#),
      2307 => to_slv(opcode_type, 16#10#),
      2308 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#03#),
      2337 => to_slv(opcode_type, 16#02#),
      2338 => to_slv(opcode_type, 16#01#),
      2339 => to_slv(opcode_type, 16#5E#),
      2340 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#05#),
      2369 => to_slv(opcode_type, 16#04#),
      2370 => to_slv(opcode_type, 16#03#),
      2371 => to_slv(opcode_type, 16#0E#),
      2372 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#02#),
      2402 => to_slv(opcode_type, 16#0C#),
      2403 => to_slv(opcode_type, 16#0A#),
      2404 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#09#),
      2433 => to_slv(opcode_type, 16#05#),
      2434 => to_slv(opcode_type, 16#0C#),
      2435 => to_slv(opcode_type, 16#0D#),
      2436 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#05#),
      2465 => to_slv(opcode_type, 16#05#),
      2466 => to_slv(opcode_type, 16#04#),
      2467 => to_slv(opcode_type, 16#0F#),
      2468 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#05#),
      2497 => to_slv(opcode_type, 16#07#),
      2498 => to_slv(opcode_type, 16#0D#),
      2499 => to_slv(opcode_type, 16#11#),
      2500 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#09#),
      2529 => to_slv(opcode_type, 16#05#),
      2530 => to_slv(opcode_type, 16#11#),
      2531 => to_slv(opcode_type, 16#0C#),
      2532 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#07#),
      2561 => to_slv(opcode_type, 16#04#),
      2562 => to_slv(opcode_type, 16#10#),
      2563 => to_slv(opcode_type, 16#0B#),
      2564 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#07#),
      2593 => to_slv(opcode_type, 16#05#),
      2594 => to_slv(opcode_type, 16#0D#),
      2595 => to_slv(opcode_type, 16#10#),
      2596 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#08#),
      2625 => to_slv(opcode_type, 16#01#),
      2626 => to_slv(opcode_type, 16#0C#),
      2627 => to_slv(opcode_type, 16#80#),
      2628 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#03#),
      2657 => to_slv(opcode_type, 16#05#),
      2658 => to_slv(opcode_type, 16#02#),
      2659 => to_slv(opcode_type, 16#0A#),
      2660 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#05#),
      2689 => to_slv(opcode_type, 16#07#),
      2690 => to_slv(opcode_type, 16#0B#),
      2691 => to_slv(opcode_type, 16#0D#),
      2692 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#09#),
      2721 => to_slv(opcode_type, 16#01#),
      2722 => to_slv(opcode_type, 16#0E#),
      2723 => to_slv(opcode_type, 16#11#),
      2724 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#07#),
      2753 => to_slv(opcode_type, 16#05#),
      2754 => to_slv(opcode_type, 16#10#),
      2755 => to_slv(opcode_type, 16#10#),
      2756 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#05#),
      2785 => to_slv(opcode_type, 16#07#),
      2786 => to_slv(opcode_type, 16#0D#),
      2787 => to_slv(opcode_type, 16#0A#),
      2788 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#08#),
      2817 => to_slv(opcode_type, 16#05#),
      2818 => to_slv(opcode_type, 16#0B#),
      2819 => to_slv(opcode_type, 16#0A#),
      2820 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#09#),
      2849 => to_slv(opcode_type, 16#04#),
      2850 => to_slv(opcode_type, 16#0D#),
      2851 => to_slv(opcode_type, 16#11#),
      2852 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#02#),
      2881 => to_slv(opcode_type, 16#04#),
      2882 => to_slv(opcode_type, 16#05#),
      2883 => to_slv(opcode_type, 16#0F#),
      2884 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#02#),
      2913 => to_slv(opcode_type, 16#08#),
      2914 => to_slv(opcode_type, 16#11#),
      2915 => to_slv(opcode_type, 16#11#),
      2916 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#03#),
      2945 => to_slv(opcode_type, 16#04#),
      2946 => to_slv(opcode_type, 16#03#),
      2947 => to_slv(opcode_type, 16#0F#),
      2948 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#01#),
      2977 => to_slv(opcode_type, 16#09#),
      2978 => to_slv(opcode_type, 16#0A#),
      2979 => to_slv(opcode_type, 16#0E#),
      2980 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#07#),
      3009 => to_slv(opcode_type, 16#02#),
      3010 => to_slv(opcode_type, 16#0A#),
      3011 => to_slv(opcode_type, 16#0B#),
      3012 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#09#),
      3041 => to_slv(opcode_type, 16#04#),
      3042 => to_slv(opcode_type, 16#0B#),
      3043 => to_slv(opcode_type, 16#0F#),
      3044 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#09#),
      3073 => to_slv(opcode_type, 16#05#),
      3074 => to_slv(opcode_type, 16#0A#),
      3075 => to_slv(opcode_type, 16#0B#),
      3076 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#07#),
      3105 => to_slv(opcode_type, 16#01#),
      3106 => to_slv(opcode_type, 16#0D#),
      3107 => to_slv(opcode_type, 16#0B#),
      3108 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#08#),
      3137 => to_slv(opcode_type, 16#01#),
      3138 => to_slv(opcode_type, 16#0A#),
      3139 => to_slv(opcode_type, 16#0D#),
      3140 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#01#),
      3169 => to_slv(opcode_type, 16#06#),
      3170 => to_slv(opcode_type, 16#BD#),
      3171 => to_slv(opcode_type, 16#11#),
      3172 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#07#),
      3201 => to_slv(opcode_type, 16#04#),
      3202 => to_slv(opcode_type, 16#0E#),
      3203 => to_slv(opcode_type, 16#11#),
      3204 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#01#),
      3233 => to_slv(opcode_type, 16#08#),
      3234 => to_slv(opcode_type, 16#11#),
      3235 => to_slv(opcode_type, 16#0F#),
      3236 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#09#),
      3265 => to_slv(opcode_type, 16#04#),
      3266 => to_slv(opcode_type, 16#0D#),
      3267 => to_slv(opcode_type, 16#BD#),
      3268 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#09#),
      3297 => to_slv(opcode_type, 16#01#),
      3298 => to_slv(opcode_type, 16#10#),
      3299 => to_slv(opcode_type, 16#10#),
      3300 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#08#),
      3329 => to_slv(opcode_type, 16#04#),
      3330 => to_slv(opcode_type, 16#0F#),
      3331 => to_slv(opcode_type, 16#0D#),
      3332 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#03#),
      3361 => to_slv(opcode_type, 16#03#),
      3362 => to_slv(opcode_type, 16#04#),
      3363 => to_slv(opcode_type, 16#CA#),
      3364 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#02#),
      3393 => to_slv(opcode_type, 16#01#),
      3394 => to_slv(opcode_type, 16#01#),
      3395 => to_slv(opcode_type, 16#0A#),
      3396 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#07#),
      3425 => to_slv(opcode_type, 16#01#),
      3426 => to_slv(opcode_type, 16#11#),
      3427 => to_slv(opcode_type, 16#0C#),
      3428 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#03#),
      3457 => to_slv(opcode_type, 16#03#),
      3458 => to_slv(opcode_type, 16#04#),
      3459 => to_slv(opcode_type, 16#0A#),
      3460 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#03#),
      3489 => to_slv(opcode_type, 16#06#),
      3490 => to_slv(opcode_type, 16#0C#),
      3491 => to_slv(opcode_type, 16#0C#),
      3492 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#08#),
      3521 => to_slv(opcode_type, 16#02#),
      3522 => to_slv(opcode_type, 16#0D#),
      3523 => to_slv(opcode_type, 16#0F#),
      3524 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#03#),
      3553 => to_slv(opcode_type, 16#08#),
      3554 => to_slv(opcode_type, 16#0B#),
      3555 => to_slv(opcode_type, 16#0E#),
      3556 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#01#),
      3585 => to_slv(opcode_type, 16#03#),
      3586 => to_slv(opcode_type, 16#01#),
      3587 => to_slv(opcode_type, 16#0C#),
      3588 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#09#),
      3617 => to_slv(opcode_type, 16#02#),
      3618 => to_slv(opcode_type, 16#0A#),
      3619 => to_slv(opcode_type, 16#10#),
      3620 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#06#),
      3649 => to_slv(opcode_type, 16#03#),
      3650 => to_slv(opcode_type, 16#0E#),
      3651 => to_slv(opcode_type, 16#0D#),
      3652 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#04#),
      3681 => to_slv(opcode_type, 16#05#),
      3682 => to_slv(opcode_type, 16#04#),
      3683 => to_slv(opcode_type, 16#0B#),
      3684 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#09#),
      3713 => to_slv(opcode_type, 16#04#),
      3714 => to_slv(opcode_type, 16#0E#),
      3715 => to_slv(opcode_type, 16#10#),
      3716 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#06#),
      3745 => to_slv(opcode_type, 16#02#),
      3746 => to_slv(opcode_type, 16#0D#),
      3747 => to_slv(opcode_type, 16#0C#),
      3748 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#05#),
      3777 => to_slv(opcode_type, 16#02#),
      3778 => to_slv(opcode_type, 16#03#),
      3779 => to_slv(opcode_type, 16#C6#),
      3780 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#05#),
      3809 => to_slv(opcode_type, 16#03#),
      3810 => to_slv(opcode_type, 16#03#),
      3811 => to_slv(opcode_type, 16#10#),
      3812 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#09#),
      3841 => to_slv(opcode_type, 16#03#),
      3842 => to_slv(opcode_type, 16#11#),
      3843 => to_slv(opcode_type, 16#0D#),
      3844 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#01#),
      3873 => to_slv(opcode_type, 16#03#),
      3874 => to_slv(opcode_type, 16#05#),
      3875 => to_slv(opcode_type, 16#10#),
      3876 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#04#),
      3905 => to_slv(opcode_type, 16#03#),
      3906 => to_slv(opcode_type, 16#04#),
      3907 => to_slv(opcode_type, 16#0F#),
      3908 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#05#),
      3937 => to_slv(opcode_type, 16#06#),
      3938 => to_slv(opcode_type, 16#F3#),
      3939 => to_slv(opcode_type, 16#0C#),
      3940 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#01#),
      3969 => to_slv(opcode_type, 16#02#),
      3970 => to_slv(opcode_type, 16#04#),
      3971 => to_slv(opcode_type, 16#0C#),
      3972 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#09#),
      4001 => to_slv(opcode_type, 16#04#),
      4002 => to_slv(opcode_type, 16#0E#),
      4003 => to_slv(opcode_type, 16#0F#),
      4004 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#07#),
      4033 => to_slv(opcode_type, 16#03#),
      4034 => to_slv(opcode_type, 16#0E#),
      4035 => to_slv(opcode_type, 16#10#),
      4036 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#01#),
      4065 => to_slv(opcode_type, 16#03#),
      4066 => to_slv(opcode_type, 16#02#),
      4067 => to_slv(opcode_type, 16#0F#),
      4068 to 4095 => (others => '0')
  ),

    -- Bin `5`...
    4 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#06#),
      1 => to_slv(opcode_type, 16#06#),
      2 => to_slv(opcode_type, 16#0E#),
      3 => to_slv(opcode_type, 16#0B#),
      4 => to_slv(opcode_type, 16#0B#),
      5 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#03#),
      33 => to_slv(opcode_type, 16#06#),
      34 => to_slv(opcode_type, 16#04#),
      35 => to_slv(opcode_type, 16#0C#),
      36 => to_slv(opcode_type, 16#10#),
      37 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#02#),
      65 => to_slv(opcode_type, 16#01#),
      66 => to_slv(opcode_type, 16#08#),
      67 => to_slv(opcode_type, 16#0E#),
      68 => to_slv(opcode_type, 16#0D#),
      69 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#08#),
      97 => to_slv(opcode_type, 16#07#),
      98 => to_slv(opcode_type, 16#0F#),
      99 => to_slv(opcode_type, 16#0D#),
      100 => to_slv(opcode_type, 16#0B#),
      101 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#04#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#05#),
      131 => to_slv(opcode_type, 16#11#),
      132 => to_slv(opcode_type, 16#0D#),
      133 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#05#),
      161 => to_slv(opcode_type, 16#04#),
      162 => to_slv(opcode_type, 16#04#),
      163 => to_slv(opcode_type, 16#01#),
      164 => to_slv(opcode_type, 16#0A#),
      165 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#08#),
      193 => to_slv(opcode_type, 16#06#),
      194 => to_slv(opcode_type, 16#11#),
      195 => to_slv(opcode_type, 16#0A#),
      196 => to_slv(opcode_type, 16#0E#),
      197 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#04#),
      225 => to_slv(opcode_type, 16#07#),
      226 => to_slv(opcode_type, 16#01#),
      227 => to_slv(opcode_type, 16#10#),
      228 => to_slv(opcode_type, 16#11#),
      229 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#03#),
      257 => to_slv(opcode_type, 16#06#),
      258 => to_slv(opcode_type, 16#04#),
      259 => to_slv(opcode_type, 16#0E#),
      260 => to_slv(opcode_type, 16#0E#),
      261 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#03#),
      289 => to_slv(opcode_type, 16#08#),
      290 => to_slv(opcode_type, 16#02#),
      291 => to_slv(opcode_type, 16#0C#),
      292 => to_slv(opcode_type, 16#10#),
      293 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#07#),
      321 => to_slv(opcode_type, 16#08#),
      322 => to_slv(opcode_type, 16#0B#),
      323 => to_slv(opcode_type, 16#0E#),
      324 => to_slv(opcode_type, 16#0E#),
      325 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#09#),
      353 => to_slv(opcode_type, 16#08#),
      354 => to_slv(opcode_type, 16#93#),
      355 => to_slv(opcode_type, 16#0E#),
      356 => to_slv(opcode_type, 16#0E#),
      357 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#06#),
      385 => to_slv(opcode_type, 16#09#),
      386 => to_slv(opcode_type, 16#0F#),
      387 => to_slv(opcode_type, 16#0C#),
      388 => to_slv(opcode_type, 16#0E#),
      389 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#06#),
      417 => to_slv(opcode_type, 16#06#),
      418 => to_slv(opcode_type, 16#11#),
      419 => to_slv(opcode_type, 16#0A#),
      420 => to_slv(opcode_type, 16#0B#),
      421 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#09#),
      449 => to_slv(opcode_type, 16#03#),
      450 => to_slv(opcode_type, 16#01#),
      451 => to_slv(opcode_type, 16#10#),
      452 => to_slv(opcode_type, 16#0D#),
      453 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#04#),
      481 => to_slv(opcode_type, 16#05#),
      482 => to_slv(opcode_type, 16#09#),
      483 => to_slv(opcode_type, 16#11#),
      484 => to_slv(opcode_type, 16#0E#),
      485 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#03#),
      514 => to_slv(opcode_type, 16#04#),
      515 => to_slv(opcode_type, 16#0C#),
      516 => to_slv(opcode_type, 16#11#),
      517 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#05#),
      545 => to_slv(opcode_type, 16#02#),
      546 => to_slv(opcode_type, 16#05#),
      547 => to_slv(opcode_type, 16#02#),
      548 => to_slv(opcode_type, 16#11#),
      549 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#02#),
      577 => to_slv(opcode_type, 16#06#),
      578 => to_slv(opcode_type, 16#03#),
      579 => to_slv(opcode_type, 16#11#),
      580 => to_slv(opcode_type, 16#0C#),
      581 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#01#),
      609 => to_slv(opcode_type, 16#04#),
      610 => to_slv(opcode_type, 16#01#),
      611 => to_slv(opcode_type, 16#05#),
      612 => to_slv(opcode_type, 16#11#),
      613 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#01#),
      641 => to_slv(opcode_type, 16#01#),
      642 => to_slv(opcode_type, 16#07#),
      643 => to_slv(opcode_type, 16#0D#),
      644 => to_slv(opcode_type, 16#FE#),
      645 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#08#),
      673 => to_slv(opcode_type, 16#04#),
      674 => to_slv(opcode_type, 16#05#),
      675 => to_slv(opcode_type, 16#0C#),
      676 => to_slv(opcode_type, 16#0F#),
      677 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#04#),
      705 => to_slv(opcode_type, 16#07#),
      706 => to_slv(opcode_type, 16#03#),
      707 => to_slv(opcode_type, 16#0F#),
      708 => to_slv(opcode_type, 16#11#),
      709 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#03#),
      737 => to_slv(opcode_type, 16#07#),
      738 => to_slv(opcode_type, 16#02#),
      739 => to_slv(opcode_type, 16#0C#),
      740 => to_slv(opcode_type, 16#0F#),
      741 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#04#),
      769 => to_slv(opcode_type, 16#04#),
      770 => to_slv(opcode_type, 16#01#),
      771 => to_slv(opcode_type, 16#02#),
      772 => to_slv(opcode_type, 16#0D#),
      773 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#02#),
      801 => to_slv(opcode_type, 16#03#),
      802 => to_slv(opcode_type, 16#03#),
      803 => to_slv(opcode_type, 16#04#),
      804 => to_slv(opcode_type, 16#0D#),
      805 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#02#),
      833 => to_slv(opcode_type, 16#01#),
      834 => to_slv(opcode_type, 16#09#),
      835 => to_slv(opcode_type, 16#0C#),
      836 => to_slv(opcode_type, 16#0C#),
      837 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#06#),
      865 => to_slv(opcode_type, 16#08#),
      866 => to_slv(opcode_type, 16#11#),
      867 => to_slv(opcode_type, 16#10#),
      868 => to_slv(opcode_type, 16#0C#),
      869 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#03#),
      897 => to_slv(opcode_type, 16#07#),
      898 => to_slv(opcode_type, 16#04#),
      899 => to_slv(opcode_type, 16#10#),
      900 => to_slv(opcode_type, 16#0A#),
      901 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#02#),
      929 => to_slv(opcode_type, 16#06#),
      930 => to_slv(opcode_type, 16#05#),
      931 => to_slv(opcode_type, 16#0D#),
      932 => to_slv(opcode_type, 16#0A#),
      933 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#03#),
      961 => to_slv(opcode_type, 16#05#),
      962 => to_slv(opcode_type, 16#09#),
      963 => to_slv(opcode_type, 16#0F#),
      964 => to_slv(opcode_type, 16#10#),
      965 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#09#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#0C#),
      995 => to_slv(opcode_type, 16#0B#),
      996 => to_slv(opcode_type, 16#0F#),
      997 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#04#),
      1025 => to_slv(opcode_type, 16#04#),
      1026 => to_slv(opcode_type, 16#09#),
      1027 => to_slv(opcode_type, 16#0B#),
      1028 => to_slv(opcode_type, 16#0A#),
      1029 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#07#),
      1057 => to_slv(opcode_type, 16#06#),
      1058 => to_slv(opcode_type, 16#10#),
      1059 => to_slv(opcode_type, 16#0E#),
      1060 => to_slv(opcode_type, 16#0B#),
      1061 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#08#),
      1089 => to_slv(opcode_type, 16#09#),
      1090 => to_slv(opcode_type, 16#0D#),
      1091 => to_slv(opcode_type, 16#0F#),
      1092 => to_slv(opcode_type, 16#0D#),
      1093 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#06#),
      1121 => to_slv(opcode_type, 16#04#),
      1122 => to_slv(opcode_type, 16#05#),
      1123 => to_slv(opcode_type, 16#0D#),
      1124 => to_slv(opcode_type, 16#EC#),
      1125 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#05#),
      1153 => to_slv(opcode_type, 16#01#),
      1154 => to_slv(opcode_type, 16#05#),
      1155 => to_slv(opcode_type, 16#03#),
      1156 => to_slv(opcode_type, 16#0B#),
      1157 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#09#),
      1185 => to_slv(opcode_type, 16#05#),
      1186 => to_slv(opcode_type, 16#05#),
      1187 => to_slv(opcode_type, 16#10#),
      1188 => to_slv(opcode_type, 16#0F#),
      1189 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#07#),
      1217 => to_slv(opcode_type, 16#06#),
      1218 => to_slv(opcode_type, 16#10#),
      1219 => to_slv(opcode_type, 16#0E#),
      1220 => to_slv(opcode_type, 16#0A#),
      1221 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#05#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#01#),
      1251 => to_slv(opcode_type, 16#0F#),
      1252 => to_slv(opcode_type, 16#11#),
      1253 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#07#),
      1281 => to_slv(opcode_type, 16#04#),
      1282 => to_slv(opcode_type, 16#01#),
      1283 => to_slv(opcode_type, 16#0F#),
      1284 => to_slv(opcode_type, 16#0E#),
      1285 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#03#),
      1313 => to_slv(opcode_type, 16#06#),
      1314 => to_slv(opcode_type, 16#04#),
      1315 => to_slv(opcode_type, 16#0F#),
      1316 => to_slv(opcode_type, 16#99#),
      1317 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#06#),
      1345 => to_slv(opcode_type, 16#08#),
      1346 => to_slv(opcode_type, 16#0D#),
      1347 => to_slv(opcode_type, 16#C4#),
      1348 => to_slv(opcode_type, 16#0E#),
      1349 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#07#),
      1377 => to_slv(opcode_type, 16#03#),
      1378 => to_slv(opcode_type, 16#01#),
      1379 => to_slv(opcode_type, 16#34#),
      1380 => to_slv(opcode_type, 16#0E#),
      1381 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#09#),
      1409 => to_slv(opcode_type, 16#02#),
      1410 => to_slv(opcode_type, 16#04#),
      1411 => to_slv(opcode_type, 16#0F#),
      1412 => to_slv(opcode_type, 16#0F#),
      1413 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#09#),
      1441 => to_slv(opcode_type, 16#09#),
      1442 => to_slv(opcode_type, 16#0C#),
      1443 => to_slv(opcode_type, 16#0E#),
      1444 => to_slv(opcode_type, 16#11#),
      1445 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#02#),
      1473 => to_slv(opcode_type, 16#01#),
      1474 => to_slv(opcode_type, 16#02#),
      1475 => to_slv(opcode_type, 16#01#),
      1476 => to_slv(opcode_type, 16#0E#),
      1477 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#08#),
      1505 => to_slv(opcode_type, 16#07#),
      1506 => to_slv(opcode_type, 16#0A#),
      1507 => to_slv(opcode_type, 16#10#),
      1508 => to_slv(opcode_type, 16#0D#),
      1509 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#05#),
      1537 => to_slv(opcode_type, 16#09#),
      1538 => to_slv(opcode_type, 16#03#),
      1539 => to_slv(opcode_type, 16#88#),
      1540 => to_slv(opcode_type, 16#10#),
      1541 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#05#),
      1569 => to_slv(opcode_type, 16#04#),
      1570 => to_slv(opcode_type, 16#04#),
      1571 => to_slv(opcode_type, 16#02#),
      1572 => to_slv(opcode_type, 16#0E#),
      1573 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#08#),
      1601 => to_slv(opcode_type, 16#08#),
      1602 => to_slv(opcode_type, 16#0C#),
      1603 => to_slv(opcode_type, 16#10#),
      1604 => to_slv(opcode_type, 16#0C#),
      1605 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#05#),
      1633 => to_slv(opcode_type, 16#02#),
      1634 => to_slv(opcode_type, 16#02#),
      1635 => to_slv(opcode_type, 16#04#),
      1636 => to_slv(opcode_type, 16#10#),
      1637 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#02#),
      1665 => to_slv(opcode_type, 16#03#),
      1666 => to_slv(opcode_type, 16#03#),
      1667 => to_slv(opcode_type, 16#05#),
      1668 => to_slv(opcode_type, 16#0A#),
      1669 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#04#),
      1697 => to_slv(opcode_type, 16#05#),
      1698 => to_slv(opcode_type, 16#07#),
      1699 => to_slv(opcode_type, 16#0A#),
      1700 => to_slv(opcode_type, 16#0B#),
      1701 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#04#),
      1729 => to_slv(opcode_type, 16#09#),
      1730 => to_slv(opcode_type, 16#02#),
      1731 => to_slv(opcode_type, 16#0C#),
      1732 => to_slv(opcode_type, 16#0D#),
      1733 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#02#),
      1761 => to_slv(opcode_type, 16#01#),
      1762 => to_slv(opcode_type, 16#01#),
      1763 => to_slv(opcode_type, 16#02#),
      1764 => to_slv(opcode_type, 16#41#),
      1765 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#09#),
      1793 => to_slv(opcode_type, 16#05#),
      1794 => to_slv(opcode_type, 16#01#),
      1795 => to_slv(opcode_type, 16#0B#),
      1796 => to_slv(opcode_type, 16#11#),
      1797 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#06#),
      1825 => to_slv(opcode_type, 16#04#),
      1826 => to_slv(opcode_type, 16#02#),
      1827 => to_slv(opcode_type, 16#0B#),
      1828 => to_slv(opcode_type, 16#2B#),
      1829 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#01#),
      1857 => to_slv(opcode_type, 16#08#),
      1858 => to_slv(opcode_type, 16#05#),
      1859 => to_slv(opcode_type, 16#0C#),
      1860 => to_slv(opcode_type, 16#0F#),
      1861 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#03#),
      1889 => to_slv(opcode_type, 16#04#),
      1890 => to_slv(opcode_type, 16#06#),
      1891 => to_slv(opcode_type, 16#0C#),
      1892 => to_slv(opcode_type, 16#0F#),
      1893 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#02#),
      1921 => to_slv(opcode_type, 16#02#),
      1922 => to_slv(opcode_type, 16#02#),
      1923 => to_slv(opcode_type, 16#05#),
      1924 => to_slv(opcode_type, 16#0C#),
      1925 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#03#),
      1953 => to_slv(opcode_type, 16#01#),
      1954 => to_slv(opcode_type, 16#01#),
      1955 => to_slv(opcode_type, 16#01#),
      1956 => to_slv(opcode_type, 16#2E#),
      1957 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#05#),
      1985 => to_slv(opcode_type, 16#04#),
      1986 => to_slv(opcode_type, 16#02#),
      1987 => to_slv(opcode_type, 16#03#),
      1988 => to_slv(opcode_type, 16#0A#),
      1989 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#04#),
      2017 => to_slv(opcode_type, 16#02#),
      2018 => to_slv(opcode_type, 16#07#),
      2019 => to_slv(opcode_type, 16#0D#),
      2020 => to_slv(opcode_type, 16#0D#),
      2021 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#07#),
      2049 => to_slv(opcode_type, 16#06#),
      2050 => to_slv(opcode_type, 16#11#),
      2051 => to_slv(opcode_type, 16#0A#),
      2052 => to_slv(opcode_type, 16#C6#),
      2053 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#07#),
      2081 => to_slv(opcode_type, 16#07#),
      2082 => to_slv(opcode_type, 16#0D#),
      2083 => to_slv(opcode_type, 16#0C#),
      2084 => to_slv(opcode_type, 16#11#),
      2085 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#05#),
      2113 => to_slv(opcode_type, 16#04#),
      2114 => to_slv(opcode_type, 16#03#),
      2115 => to_slv(opcode_type, 16#04#),
      2116 => to_slv(opcode_type, 16#0F#),
      2117 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#06#),
      2145 => to_slv(opcode_type, 16#09#),
      2146 => to_slv(opcode_type, 16#0C#),
      2147 => to_slv(opcode_type, 16#0B#),
      2148 => to_slv(opcode_type, 16#0D#),
      2149 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#05#),
      2177 => to_slv(opcode_type, 16#02#),
      2178 => to_slv(opcode_type, 16#01#),
      2179 => to_slv(opcode_type, 16#04#),
      2180 => to_slv(opcode_type, 16#10#),
      2181 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#05#),
      2209 => to_slv(opcode_type, 16#01#),
      2210 => to_slv(opcode_type, 16#09#),
      2211 => to_slv(opcode_type, 16#0A#),
      2212 => to_slv(opcode_type, 16#1F#),
      2213 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#06#),
      2242 => to_slv(opcode_type, 16#0A#),
      2243 => to_slv(opcode_type, 16#0B#),
      2244 => to_slv(opcode_type, 16#0E#),
      2245 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#08#),
      2273 => to_slv(opcode_type, 16#03#),
      2274 => to_slv(opcode_type, 16#03#),
      2275 => to_slv(opcode_type, 16#11#),
      2276 => to_slv(opcode_type, 16#0C#),
      2277 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#02#),
      2305 => to_slv(opcode_type, 16#04#),
      2306 => to_slv(opcode_type, 16#03#),
      2307 => to_slv(opcode_type, 16#03#),
      2308 => to_slv(opcode_type, 16#34#),
      2309 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#01#),
      2337 => to_slv(opcode_type, 16#03#),
      2338 => to_slv(opcode_type, 16#05#),
      2339 => to_slv(opcode_type, 16#05#),
      2340 => to_slv(opcode_type, 16#0A#),
      2341 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#02#),
      2369 => to_slv(opcode_type, 16#07#),
      2370 => to_slv(opcode_type, 16#03#),
      2371 => to_slv(opcode_type, 16#0D#),
      2372 => to_slv(opcode_type, 16#0A#),
      2373 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#09#),
      2401 => to_slv(opcode_type, 16#02#),
      2402 => to_slv(opcode_type, 16#01#),
      2403 => to_slv(opcode_type, 16#B7#),
      2404 => to_slv(opcode_type, 16#11#),
      2405 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#01#),
      2433 => to_slv(opcode_type, 16#03#),
      2434 => to_slv(opcode_type, 16#09#),
      2435 => to_slv(opcode_type, 16#11#),
      2436 => to_slv(opcode_type, 16#0C#),
      2437 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#04#),
      2465 => to_slv(opcode_type, 16#04#),
      2466 => to_slv(opcode_type, 16#07#),
      2467 => to_slv(opcode_type, 16#0C#),
      2468 => to_slv(opcode_type, 16#10#),
      2469 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#05#),
      2497 => to_slv(opcode_type, 16#02#),
      2498 => to_slv(opcode_type, 16#07#),
      2499 => to_slv(opcode_type, 16#0F#),
      2500 => to_slv(opcode_type, 16#0D#),
      2501 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#03#),
      2529 => to_slv(opcode_type, 16#07#),
      2530 => to_slv(opcode_type, 16#01#),
      2531 => to_slv(opcode_type, 16#0C#),
      2532 => to_slv(opcode_type, 16#0D#),
      2533 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#04#),
      2561 => to_slv(opcode_type, 16#08#),
      2562 => to_slv(opcode_type, 16#05#),
      2563 => to_slv(opcode_type, 16#0C#),
      2564 => to_slv(opcode_type, 16#11#),
      2565 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#08#),
      2593 => to_slv(opcode_type, 16#06#),
      2594 => to_slv(opcode_type, 16#E0#),
      2595 => to_slv(opcode_type, 16#11#),
      2596 => to_slv(opcode_type, 16#0B#),
      2597 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#02#),
      2625 => to_slv(opcode_type, 16#04#),
      2626 => to_slv(opcode_type, 16#04#),
      2627 => to_slv(opcode_type, 16#04#),
      2628 => to_slv(opcode_type, 16#10#),
      2629 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#07#),
      2657 => to_slv(opcode_type, 16#03#),
      2658 => to_slv(opcode_type, 16#03#),
      2659 => to_slv(opcode_type, 16#0D#),
      2660 => to_slv(opcode_type, 16#0E#),
      2661 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#06#),
      2689 => to_slv(opcode_type, 16#05#),
      2690 => to_slv(opcode_type, 16#03#),
      2691 => to_slv(opcode_type, 16#10#),
      2692 => to_slv(opcode_type, 16#0E#),
      2693 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#08#),
      2721 => to_slv(opcode_type, 16#02#),
      2722 => to_slv(opcode_type, 16#04#),
      2723 => to_slv(opcode_type, 16#0E#),
      2724 => to_slv(opcode_type, 16#0A#),
      2725 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#03#),
      2753 => to_slv(opcode_type, 16#04#),
      2754 => to_slv(opcode_type, 16#09#),
      2755 => to_slv(opcode_type, 16#0F#),
      2756 => to_slv(opcode_type, 16#0F#),
      2757 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#03#),
      2785 => to_slv(opcode_type, 16#09#),
      2786 => to_slv(opcode_type, 16#03#),
      2787 => to_slv(opcode_type, 16#11#),
      2788 => to_slv(opcode_type, 16#0B#),
      2789 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#07#),
      2817 => to_slv(opcode_type, 16#04#),
      2818 => to_slv(opcode_type, 16#05#),
      2819 => to_slv(opcode_type, 16#0D#),
      2820 => to_slv(opcode_type, 16#11#),
      2821 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#01#),
      2849 => to_slv(opcode_type, 16#08#),
      2850 => to_slv(opcode_type, 16#05#),
      2851 => to_slv(opcode_type, 16#0D#),
      2852 => to_slv(opcode_type, 16#0C#),
      2853 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#09#),
      2881 => to_slv(opcode_type, 16#01#),
      2882 => to_slv(opcode_type, 16#05#),
      2883 => to_slv(opcode_type, 16#0E#),
      2884 => to_slv(opcode_type, 16#0D#),
      2885 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#02#),
      2913 => to_slv(opcode_type, 16#07#),
      2914 => to_slv(opcode_type, 16#02#),
      2915 => to_slv(opcode_type, 16#11#),
      2916 => to_slv(opcode_type, 16#0B#),
      2917 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#06#),
      2945 => to_slv(opcode_type, 16#01#),
      2946 => to_slv(opcode_type, 16#04#),
      2947 => to_slv(opcode_type, 16#10#),
      2948 => to_slv(opcode_type, 16#0B#),
      2949 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#09#),
      2977 => to_slv(opcode_type, 16#07#),
      2978 => to_slv(opcode_type, 16#0B#),
      2979 => to_slv(opcode_type, 16#10#),
      2980 => to_slv(opcode_type, 16#0F#),
      2981 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#02#),
      3009 => to_slv(opcode_type, 16#05#),
      3010 => to_slv(opcode_type, 16#08#),
      3011 => to_slv(opcode_type, 16#0D#),
      3012 => to_slv(opcode_type, 16#0E#),
      3013 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#01#),
      3041 => to_slv(opcode_type, 16#03#),
      3042 => to_slv(opcode_type, 16#08#),
      3043 => to_slv(opcode_type, 16#0A#),
      3044 => to_slv(opcode_type, 16#0F#),
      3045 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#03#),
      3073 => to_slv(opcode_type, 16#09#),
      3074 => to_slv(opcode_type, 16#03#),
      3075 => to_slv(opcode_type, 16#11#),
      3076 => to_slv(opcode_type, 16#0C#),
      3077 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#06#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#11#),
      3107 => to_slv(opcode_type, 16#0D#),
      3108 => to_slv(opcode_type, 16#15#),
      3109 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#08#),
      3137 => to_slv(opcode_type, 16#01#),
      3138 => to_slv(opcode_type, 16#03#),
      3139 => to_slv(opcode_type, 16#0F#),
      3140 => to_slv(opcode_type, 16#11#),
      3141 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#03#),
      3169 => to_slv(opcode_type, 16#02#),
      3170 => to_slv(opcode_type, 16#08#),
      3171 => to_slv(opcode_type, 16#0F#),
      3172 => to_slv(opcode_type, 16#E1#),
      3173 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#03#),
      3201 => to_slv(opcode_type, 16#08#),
      3202 => to_slv(opcode_type, 16#04#),
      3203 => to_slv(opcode_type, 16#0B#),
      3204 => to_slv(opcode_type, 16#0C#),
      3205 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#05#),
      3233 => to_slv(opcode_type, 16#08#),
      3234 => to_slv(opcode_type, 16#05#),
      3235 => to_slv(opcode_type, 16#0A#),
      3236 => to_slv(opcode_type, 16#0C#),
      3237 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#08#),
      3265 => to_slv(opcode_type, 16#02#),
      3266 => to_slv(opcode_type, 16#04#),
      3267 => to_slv(opcode_type, 16#FB#),
      3268 => to_slv(opcode_type, 16#0E#),
      3269 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#08#),
      3297 => to_slv(opcode_type, 16#03#),
      3298 => to_slv(opcode_type, 16#05#),
      3299 => to_slv(opcode_type, 16#63#),
      3300 => to_slv(opcode_type, 16#86#),
      3301 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#01#),
      3329 => to_slv(opcode_type, 16#02#),
      3330 => to_slv(opcode_type, 16#08#),
      3331 => to_slv(opcode_type, 16#6F#),
      3332 => to_slv(opcode_type, 16#0F#),
      3333 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#01#),
      3361 => to_slv(opcode_type, 16#02#),
      3362 => to_slv(opcode_type, 16#06#),
      3363 => to_slv(opcode_type, 16#0B#),
      3364 => to_slv(opcode_type, 16#0A#),
      3365 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#09#),
      3393 => to_slv(opcode_type, 16#09#),
      3394 => to_slv(opcode_type, 16#0F#),
      3395 => to_slv(opcode_type, 16#0E#),
      3396 => to_slv(opcode_type, 16#0B#),
      3397 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#01#),
      3425 => to_slv(opcode_type, 16#05#),
      3426 => to_slv(opcode_type, 16#05#),
      3427 => to_slv(opcode_type, 16#01#),
      3428 => to_slv(opcode_type, 16#11#),
      3429 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#06#),
      3457 => to_slv(opcode_type, 16#04#),
      3458 => to_slv(opcode_type, 16#04#),
      3459 => to_slv(opcode_type, 16#0A#),
      3460 => to_slv(opcode_type, 16#0F#),
      3461 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#05#),
      3489 => to_slv(opcode_type, 16#03#),
      3490 => to_slv(opcode_type, 16#09#),
      3491 => to_slv(opcode_type, 16#0C#),
      3492 => to_slv(opcode_type, 16#0D#),
      3493 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#05#),
      3521 => to_slv(opcode_type, 16#03#),
      3522 => to_slv(opcode_type, 16#01#),
      3523 => to_slv(opcode_type, 16#04#),
      3524 => to_slv(opcode_type, 16#0F#),
      3525 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#09#),
      3553 => to_slv(opcode_type, 16#04#),
      3554 => to_slv(opcode_type, 16#05#),
      3555 => to_slv(opcode_type, 16#0C#),
      3556 => to_slv(opcode_type, 16#10#),
      3557 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#04#),
      3585 => to_slv(opcode_type, 16#05#),
      3586 => to_slv(opcode_type, 16#01#),
      3587 => to_slv(opcode_type, 16#01#),
      3588 => to_slv(opcode_type, 16#0C#),
      3589 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#03#),
      3617 => to_slv(opcode_type, 16#06#),
      3618 => to_slv(opcode_type, 16#04#),
      3619 => to_slv(opcode_type, 16#0E#),
      3620 => to_slv(opcode_type, 16#0D#),
      3621 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#02#),
      3649 => to_slv(opcode_type, 16#07#),
      3650 => to_slv(opcode_type, 16#04#),
      3651 => to_slv(opcode_type, 16#0E#),
      3652 => to_slv(opcode_type, 16#0F#),
      3653 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#04#),
      3681 => to_slv(opcode_type, 16#05#),
      3682 => to_slv(opcode_type, 16#05#),
      3683 => to_slv(opcode_type, 16#01#),
      3684 => to_slv(opcode_type, 16#0F#),
      3685 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#04#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#03#),
      3715 => to_slv(opcode_type, 16#73#),
      3716 => to_slv(opcode_type, 16#0A#),
      3717 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#02#),
      3745 => to_slv(opcode_type, 16#01#),
      3746 => to_slv(opcode_type, 16#03#),
      3747 => to_slv(opcode_type, 16#02#),
      3748 => to_slv(opcode_type, 16#0C#),
      3749 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#08#),
      3777 => to_slv(opcode_type, 16#07#),
      3778 => to_slv(opcode_type, 16#0B#),
      3779 => to_slv(opcode_type, 16#0F#),
      3780 => to_slv(opcode_type, 16#0B#),
      3781 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#04#),
      3809 => to_slv(opcode_type, 16#04#),
      3810 => to_slv(opcode_type, 16#02#),
      3811 => to_slv(opcode_type, 16#05#),
      3812 => to_slv(opcode_type, 16#77#),
      3813 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#02#),
      3841 => to_slv(opcode_type, 16#02#),
      3842 => to_slv(opcode_type, 16#02#),
      3843 => to_slv(opcode_type, 16#05#),
      3844 => to_slv(opcode_type, 16#0A#),
      3845 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#08#),
      3873 => to_slv(opcode_type, 16#04#),
      3874 => to_slv(opcode_type, 16#02#),
      3875 => to_slv(opcode_type, 16#BB#),
      3876 => to_slv(opcode_type, 16#0A#),
      3877 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#07#),
      3905 => to_slv(opcode_type, 16#04#),
      3906 => to_slv(opcode_type, 16#01#),
      3907 => to_slv(opcode_type, 16#CF#),
      3908 => to_slv(opcode_type, 16#A3#),
      3909 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#03#),
      3937 => to_slv(opcode_type, 16#01#),
      3938 => to_slv(opcode_type, 16#09#),
      3939 => to_slv(opcode_type, 16#0F#),
      3940 => to_slv(opcode_type, 16#0D#),
      3941 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#01#),
      3969 => to_slv(opcode_type, 16#04#),
      3970 => to_slv(opcode_type, 16#08#),
      3971 => to_slv(opcode_type, 16#0D#),
      3972 => to_slv(opcode_type, 16#0F#),
      3973 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#08#),
      4001 => to_slv(opcode_type, 16#02#),
      4002 => to_slv(opcode_type, 16#05#),
      4003 => to_slv(opcode_type, 16#73#),
      4004 => to_slv(opcode_type, 16#10#),
      4005 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#09#),
      4033 => to_slv(opcode_type, 16#02#),
      4034 => to_slv(opcode_type, 16#05#),
      4035 => to_slv(opcode_type, 16#0D#),
      4036 => to_slv(opcode_type, 16#0F#),
      4037 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#03#),
      4065 => to_slv(opcode_type, 16#07#),
      4066 => to_slv(opcode_type, 16#04#),
      4067 => to_slv(opcode_type, 16#0D#),
      4068 => to_slv(opcode_type, 16#11#),
      4069 to 4095 => (others => '0')
  ),

    -- Bin `6`...
    5 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#02#),
      1 => to_slv(opcode_type, 16#09#),
      2 => to_slv(opcode_type, 16#09#),
      3 => to_slv(opcode_type, 16#0E#),
      4 => to_slv(opcode_type, 16#0A#),
      5 => to_slv(opcode_type, 16#0B#),
      6 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#06#),
      33 => to_slv(opcode_type, 16#01#),
      34 => to_slv(opcode_type, 16#02#),
      35 => to_slv(opcode_type, 16#02#),
      36 => to_slv(opcode_type, 16#11#),
      37 => to_slv(opcode_type, 16#0E#),
      38 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#09#),
      65 => to_slv(opcode_type, 16#07#),
      66 => to_slv(opcode_type, 16#05#),
      67 => to_slv(opcode_type, 16#0B#),
      68 => to_slv(opcode_type, 16#11#),
      69 => to_slv(opcode_type, 16#0D#),
      70 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#06#),
      97 => to_slv(opcode_type, 16#01#),
      98 => to_slv(opcode_type, 16#07#),
      99 => to_slv(opcode_type, 16#11#),
      100 => to_slv(opcode_type, 16#11#),
      101 => to_slv(opcode_type, 16#0D#),
      102 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#06#),
      129 => to_slv(opcode_type, 16#06#),
      130 => to_slv(opcode_type, 16#05#),
      131 => to_slv(opcode_type, 16#0B#),
      132 => to_slv(opcode_type, 16#0D#),
      133 => to_slv(opcode_type, 16#0F#),
      134 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#05#),
      161 => to_slv(opcode_type, 16#04#),
      162 => to_slv(opcode_type, 16#07#),
      163 => to_slv(opcode_type, 16#04#),
      164 => to_slv(opcode_type, 16#0B#),
      165 => to_slv(opcode_type, 16#0F#),
      166 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#03#),
      193 => to_slv(opcode_type, 16#07#),
      194 => to_slv(opcode_type, 16#04#),
      195 => to_slv(opcode_type, 16#03#),
      196 => to_slv(opcode_type, 16#0F#),
      197 => to_slv(opcode_type, 16#0B#),
      198 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#09#),
      225 => to_slv(opcode_type, 16#01#),
      226 => to_slv(opcode_type, 16#07#),
      227 => to_slv(opcode_type, 16#0F#),
      228 => to_slv(opcode_type, 16#11#),
      229 => to_slv(opcode_type, 16#0F#),
      230 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#06#),
      257 => to_slv(opcode_type, 16#03#),
      258 => to_slv(opcode_type, 16#02#),
      259 => to_slv(opcode_type, 16#02#),
      260 => to_slv(opcode_type, 16#0C#),
      261 => to_slv(opcode_type, 16#0F#),
      262 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#01#),
      290 => to_slv(opcode_type, 16#09#),
      291 => to_slv(opcode_type, 16#0E#),
      292 => to_slv(opcode_type, 16#0B#),
      293 => to_slv(opcode_type, 16#0F#),
      294 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#06#),
      321 => to_slv(opcode_type, 16#03#),
      322 => to_slv(opcode_type, 16#08#),
      323 => to_slv(opcode_type, 16#0C#),
      324 => to_slv(opcode_type, 16#0C#),
      325 => to_slv(opcode_type, 16#0F#),
      326 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#04#),
      353 => to_slv(opcode_type, 16#06#),
      354 => to_slv(opcode_type, 16#01#),
      355 => to_slv(opcode_type, 16#03#),
      356 => to_slv(opcode_type, 16#0D#),
      357 => to_slv(opcode_type, 16#0E#),
      358 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#01#),
      385 => to_slv(opcode_type, 16#05#),
      386 => to_slv(opcode_type, 16#01#),
      387 => to_slv(opcode_type, 16#08#),
      388 => to_slv(opcode_type, 16#52#),
      389 => to_slv(opcode_type, 16#0F#),
      390 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#05#),
      417 => to_slv(opcode_type, 16#01#),
      418 => to_slv(opcode_type, 16#02#),
      419 => to_slv(opcode_type, 16#09#),
      420 => to_slv(opcode_type, 16#46#),
      421 => to_slv(opcode_type, 16#0B#),
      422 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#06#),
      449 => to_slv(opcode_type, 16#09#),
      450 => to_slv(opcode_type, 16#02#),
      451 => to_slv(opcode_type, 16#0F#),
      452 => to_slv(opcode_type, 16#0E#),
      453 => to_slv(opcode_type, 16#2A#),
      454 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#01#),
      481 => to_slv(opcode_type, 16#05#),
      482 => to_slv(opcode_type, 16#09#),
      483 => to_slv(opcode_type, 16#02#),
      484 => to_slv(opcode_type, 16#A2#),
      485 => to_slv(opcode_type, 16#0F#),
      486 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#04#),
      513 => to_slv(opcode_type, 16#04#),
      514 => to_slv(opcode_type, 16#07#),
      515 => to_slv(opcode_type, 16#02#),
      516 => to_slv(opcode_type, 16#0A#),
      517 => to_slv(opcode_type, 16#0F#),
      518 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#08#),
      545 => to_slv(opcode_type, 16#04#),
      546 => to_slv(opcode_type, 16#05#),
      547 => to_slv(opcode_type, 16#03#),
      548 => to_slv(opcode_type, 16#6A#),
      549 => to_slv(opcode_type, 16#10#),
      550 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#01#),
      577 => to_slv(opcode_type, 16#03#),
      578 => to_slv(opcode_type, 16#08#),
      579 => to_slv(opcode_type, 16#04#),
      580 => to_slv(opcode_type, 16#CB#),
      581 => to_slv(opcode_type, 16#10#),
      582 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#08#),
      609 => to_slv(opcode_type, 16#07#),
      610 => to_slv(opcode_type, 16#04#),
      611 => to_slv(opcode_type, 16#11#),
      612 => to_slv(opcode_type, 16#0E#),
      613 => to_slv(opcode_type, 16#0F#),
      614 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#02#),
      641 => to_slv(opcode_type, 16#05#),
      642 => to_slv(opcode_type, 16#09#),
      643 => to_slv(opcode_type, 16#02#),
      644 => to_slv(opcode_type, 16#F6#),
      645 => to_slv(opcode_type, 16#0E#),
      646 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#03#),
      673 => to_slv(opcode_type, 16#06#),
      674 => to_slv(opcode_type, 16#09#),
      675 => to_slv(opcode_type, 16#0D#),
      676 => to_slv(opcode_type, 16#10#),
      677 => to_slv(opcode_type, 16#11#),
      678 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#01#),
      705 => to_slv(opcode_type, 16#07#),
      706 => to_slv(opcode_type, 16#06#),
      707 => to_slv(opcode_type, 16#10#),
      708 => to_slv(opcode_type, 16#10#),
      709 => to_slv(opcode_type, 16#0E#),
      710 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#07#),
      737 => to_slv(opcode_type, 16#07#),
      738 => to_slv(opcode_type, 16#01#),
      739 => to_slv(opcode_type, 16#0D#),
      740 => to_slv(opcode_type, 16#10#),
      741 => to_slv(opcode_type, 16#0B#),
      742 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#02#),
      769 => to_slv(opcode_type, 16#02#),
      770 => to_slv(opcode_type, 16#03#),
      771 => to_slv(opcode_type, 16#07#),
      772 => to_slv(opcode_type, 16#0A#),
      773 => to_slv(opcode_type, 16#0F#),
      774 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#09#),
      801 => to_slv(opcode_type, 16#08#),
      802 => to_slv(opcode_type, 16#04#),
      803 => to_slv(opcode_type, 16#0E#),
      804 => to_slv(opcode_type, 16#0B#),
      805 => to_slv(opcode_type, 16#28#),
      806 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#08#),
      833 => to_slv(opcode_type, 16#03#),
      834 => to_slv(opcode_type, 16#06#),
      835 => to_slv(opcode_type, 16#3C#),
      836 => to_slv(opcode_type, 16#1F#),
      837 => to_slv(opcode_type, 16#0E#),
      838 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#02#),
      865 => to_slv(opcode_type, 16#03#),
      866 => to_slv(opcode_type, 16#07#),
      867 => to_slv(opcode_type, 16#04#),
      868 => to_slv(opcode_type, 16#0D#),
      869 => to_slv(opcode_type, 16#0E#),
      870 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#05#),
      897 => to_slv(opcode_type, 16#09#),
      898 => to_slv(opcode_type, 16#04#),
      899 => to_slv(opcode_type, 16#01#),
      900 => to_slv(opcode_type, 16#98#),
      901 => to_slv(opcode_type, 16#11#),
      902 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#04#),
      929 => to_slv(opcode_type, 16#07#),
      930 => to_slv(opcode_type, 16#09#),
      931 => to_slv(opcode_type, 16#0C#),
      932 => to_slv(opcode_type, 16#0B#),
      933 => to_slv(opcode_type, 16#0C#),
      934 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#06#),
      961 => to_slv(opcode_type, 16#03#),
      962 => to_slv(opcode_type, 16#01#),
      963 => to_slv(opcode_type, 16#03#),
      964 => to_slv(opcode_type, 16#52#),
      965 => to_slv(opcode_type, 16#11#),
      966 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#08#),
      993 => to_slv(opcode_type, 16#04#),
      994 => to_slv(opcode_type, 16#06#),
      995 => to_slv(opcode_type, 16#0F#),
      996 => to_slv(opcode_type, 16#11#),
      997 => to_slv(opcode_type, 16#0D#),
      998 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#03#),
      1025 => to_slv(opcode_type, 16#08#),
      1026 => to_slv(opcode_type, 16#01#),
      1027 => to_slv(opcode_type, 16#04#),
      1028 => to_slv(opcode_type, 16#0E#),
      1029 => to_slv(opcode_type, 16#0B#),
      1030 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#08#),
      1057 => to_slv(opcode_type, 16#01#),
      1058 => to_slv(opcode_type, 16#01#),
      1059 => to_slv(opcode_type, 16#03#),
      1060 => to_slv(opcode_type, 16#11#),
      1061 => to_slv(opcode_type, 16#0F#),
      1062 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#02#),
      1089 => to_slv(opcode_type, 16#09#),
      1090 => to_slv(opcode_type, 16#05#),
      1091 => to_slv(opcode_type, 16#04#),
      1092 => to_slv(opcode_type, 16#0A#),
      1093 => to_slv(opcode_type, 16#10#),
      1094 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#02#),
      1121 => to_slv(opcode_type, 16#09#),
      1122 => to_slv(opcode_type, 16#03#),
      1123 => to_slv(opcode_type, 16#02#),
      1124 => to_slv(opcode_type, 16#0E#),
      1125 => to_slv(opcode_type, 16#11#),
      1126 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#09#),
      1153 => to_slv(opcode_type, 16#02#),
      1154 => to_slv(opcode_type, 16#09#),
      1155 => to_slv(opcode_type, 16#0B#),
      1156 => to_slv(opcode_type, 16#10#),
      1157 => to_slv(opcode_type, 16#0D#),
      1158 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#01#),
      1185 => to_slv(opcode_type, 16#09#),
      1186 => to_slv(opcode_type, 16#02#),
      1187 => to_slv(opcode_type, 16#02#),
      1188 => to_slv(opcode_type, 16#0B#),
      1189 => to_slv(opcode_type, 16#0A#),
      1190 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#08#),
      1217 => to_slv(opcode_type, 16#06#),
      1218 => to_slv(opcode_type, 16#02#),
      1219 => to_slv(opcode_type, 16#0A#),
      1220 => to_slv(opcode_type, 16#0F#),
      1221 => to_slv(opcode_type, 16#0F#),
      1222 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#09#),
      1249 => to_slv(opcode_type, 16#02#),
      1250 => to_slv(opcode_type, 16#03#),
      1251 => to_slv(opcode_type, 16#03#),
      1252 => to_slv(opcode_type, 16#0B#),
      1253 => to_slv(opcode_type, 16#0D#),
      1254 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#03#),
      1281 => to_slv(opcode_type, 16#04#),
      1282 => to_slv(opcode_type, 16#06#),
      1283 => to_slv(opcode_type, 16#04#),
      1284 => to_slv(opcode_type, 16#0A#),
      1285 => to_slv(opcode_type, 16#0E#),
      1286 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#09#),
      1313 => to_slv(opcode_type, 16#03#),
      1314 => to_slv(opcode_type, 16#03#),
      1315 => to_slv(opcode_type, 16#02#),
      1316 => to_slv(opcode_type, 16#0B#),
      1317 => to_slv(opcode_type, 16#E5#),
      1318 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#04#),
      1345 => to_slv(opcode_type, 16#09#),
      1346 => to_slv(opcode_type, 16#09#),
      1347 => to_slv(opcode_type, 16#11#),
      1348 => to_slv(opcode_type, 16#0C#),
      1349 => to_slv(opcode_type, 16#0C#),
      1350 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#09#),
      1377 => to_slv(opcode_type, 16#01#),
      1378 => to_slv(opcode_type, 16#09#),
      1379 => to_slv(opcode_type, 16#0A#),
      1380 => to_slv(opcode_type, 16#0F#),
      1381 => to_slv(opcode_type, 16#0A#),
      1382 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#02#),
      1410 => to_slv(opcode_type, 16#05#),
      1411 => to_slv(opcode_type, 16#02#),
      1412 => to_slv(opcode_type, 16#11#),
      1413 => to_slv(opcode_type, 16#10#),
      1414 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#06#),
      1441 => to_slv(opcode_type, 16#07#),
      1442 => to_slv(opcode_type, 16#01#),
      1443 => to_slv(opcode_type, 16#0C#),
      1444 => to_slv(opcode_type, 16#0D#),
      1445 => to_slv(opcode_type, 16#11#),
      1446 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#04#),
      1473 => to_slv(opcode_type, 16#06#),
      1474 => to_slv(opcode_type, 16#05#),
      1475 => to_slv(opcode_type, 16#05#),
      1476 => to_slv(opcode_type, 16#0E#),
      1477 => to_slv(opcode_type, 16#3C#),
      1478 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#03#),
      1505 => to_slv(opcode_type, 16#02#),
      1506 => to_slv(opcode_type, 16#03#),
      1507 => to_slv(opcode_type, 16#09#),
      1508 => to_slv(opcode_type, 16#11#),
      1509 => to_slv(opcode_type, 16#0C#),
      1510 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#01#),
      1537 => to_slv(opcode_type, 16#01#),
      1538 => to_slv(opcode_type, 16#04#),
      1539 => to_slv(opcode_type, 16#08#),
      1540 => to_slv(opcode_type, 16#85#),
      1541 => to_slv(opcode_type, 16#0E#),
      1542 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#04#),
      1569 => to_slv(opcode_type, 16#07#),
      1570 => to_slv(opcode_type, 16#06#),
      1571 => to_slv(opcode_type, 16#0D#),
      1572 => to_slv(opcode_type, 16#0A#),
      1573 => to_slv(opcode_type, 16#0E#),
      1574 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#05#),
      1601 => to_slv(opcode_type, 16#04#),
      1602 => to_slv(opcode_type, 16#07#),
      1603 => to_slv(opcode_type, 16#03#),
      1604 => to_slv(opcode_type, 16#2A#),
      1605 => to_slv(opcode_type, 16#0B#),
      1606 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#02#),
      1633 => to_slv(opcode_type, 16#06#),
      1634 => to_slv(opcode_type, 16#05#),
      1635 => to_slv(opcode_type, 16#01#),
      1636 => to_slv(opcode_type, 16#24#),
      1637 => to_slv(opcode_type, 16#0B#),
      1638 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#07#),
      1665 => to_slv(opcode_type, 16#07#),
      1666 => to_slv(opcode_type, 16#04#),
      1667 => to_slv(opcode_type, 16#0A#),
      1668 => to_slv(opcode_type, 16#0C#),
      1669 => to_slv(opcode_type, 16#0D#),
      1670 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#02#),
      1697 => to_slv(opcode_type, 16#03#),
      1698 => to_slv(opcode_type, 16#03#),
      1699 => to_slv(opcode_type, 16#09#),
      1700 => to_slv(opcode_type, 16#0D#),
      1701 => to_slv(opcode_type, 16#0D#),
      1702 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#09#),
      1729 => to_slv(opcode_type, 16#09#),
      1730 => to_slv(opcode_type, 16#05#),
      1731 => to_slv(opcode_type, 16#10#),
      1732 => to_slv(opcode_type, 16#11#),
      1733 => to_slv(opcode_type, 16#AF#),
      1734 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#04#),
      1761 => to_slv(opcode_type, 16#07#),
      1762 => to_slv(opcode_type, 16#06#),
      1763 => to_slv(opcode_type, 16#0C#),
      1764 => to_slv(opcode_type, 16#10#),
      1765 => to_slv(opcode_type, 16#11#),
      1766 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#09#),
      1793 => to_slv(opcode_type, 16#09#),
      1794 => to_slv(opcode_type, 16#03#),
      1795 => to_slv(opcode_type, 16#0A#),
      1796 => to_slv(opcode_type, 16#0E#),
      1797 => to_slv(opcode_type, 16#0A#),
      1798 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#02#),
      1825 => to_slv(opcode_type, 16#06#),
      1826 => to_slv(opcode_type, 16#02#),
      1827 => to_slv(opcode_type, 16#03#),
      1828 => to_slv(opcode_type, 16#0A#),
      1829 => to_slv(opcode_type, 16#10#),
      1830 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#07#),
      1857 => to_slv(opcode_type, 16#09#),
      1858 => to_slv(opcode_type, 16#01#),
      1859 => to_slv(opcode_type, 16#11#),
      1860 => to_slv(opcode_type, 16#0A#),
      1861 => to_slv(opcode_type, 16#0C#),
      1862 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#02#),
      1889 => to_slv(opcode_type, 16#09#),
      1890 => to_slv(opcode_type, 16#01#),
      1891 => to_slv(opcode_type, 16#05#),
      1892 => to_slv(opcode_type, 16#10#),
      1893 => to_slv(opcode_type, 16#0B#),
      1894 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#01#),
      1921 => to_slv(opcode_type, 16#08#),
      1922 => to_slv(opcode_type, 16#01#),
      1923 => to_slv(opcode_type, 16#03#),
      1924 => to_slv(opcode_type, 16#0D#),
      1925 => to_slv(opcode_type, 16#0D#),
      1926 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#09#),
      1953 => to_slv(opcode_type, 16#06#),
      1954 => to_slv(opcode_type, 16#03#),
      1955 => to_slv(opcode_type, 16#0A#),
      1956 => to_slv(opcode_type, 16#0F#),
      1957 => to_slv(opcode_type, 16#0B#),
      1958 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#01#),
      1985 => to_slv(opcode_type, 16#08#),
      1986 => to_slv(opcode_type, 16#08#),
      1987 => to_slv(opcode_type, 16#10#),
      1988 => to_slv(opcode_type, 16#0E#),
      1989 => to_slv(opcode_type, 16#D9#),
      1990 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#02#),
      2017 => to_slv(opcode_type, 16#05#),
      2018 => to_slv(opcode_type, 16#07#),
      2019 => to_slv(opcode_type, 16#01#),
      2020 => to_slv(opcode_type, 16#0B#),
      2021 => to_slv(opcode_type, 16#0A#),
      2022 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#01#),
      2049 => to_slv(opcode_type, 16#04#),
      2050 => to_slv(opcode_type, 16#08#),
      2051 => to_slv(opcode_type, 16#02#),
      2052 => to_slv(opcode_type, 16#0B#),
      2053 => to_slv(opcode_type, 16#11#),
      2054 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#02#),
      2081 => to_slv(opcode_type, 16#05#),
      2082 => to_slv(opcode_type, 16#03#),
      2083 => to_slv(opcode_type, 16#07#),
      2084 => to_slv(opcode_type, 16#11#),
      2085 => to_slv(opcode_type, 16#11#),
      2086 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#09#),
      2113 => to_slv(opcode_type, 16#05#),
      2114 => to_slv(opcode_type, 16#01#),
      2115 => to_slv(opcode_type, 16#05#),
      2116 => to_slv(opcode_type, 16#0F#),
      2117 => to_slv(opcode_type, 16#0A#),
      2118 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#07#),
      2145 => to_slv(opcode_type, 16#05#),
      2146 => to_slv(opcode_type, 16#07#),
      2147 => to_slv(opcode_type, 16#11#),
      2148 => to_slv(opcode_type, 16#0F#),
      2149 => to_slv(opcode_type, 16#0F#),
      2150 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#05#),
      2177 => to_slv(opcode_type, 16#04#),
      2178 => to_slv(opcode_type, 16#02#),
      2179 => to_slv(opcode_type, 16#07#),
      2180 => to_slv(opcode_type, 16#99#),
      2181 => to_slv(opcode_type, 16#0E#),
      2182 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#06#),
      2209 => to_slv(opcode_type, 16#02#),
      2210 => to_slv(opcode_type, 16#04#),
      2211 => to_slv(opcode_type, 16#04#),
      2212 => to_slv(opcode_type, 16#0E#),
      2213 => to_slv(opcode_type, 16#0F#),
      2214 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#01#),
      2241 => to_slv(opcode_type, 16#02#),
      2242 => to_slv(opcode_type, 16#03#),
      2243 => to_slv(opcode_type, 16#08#),
      2244 => to_slv(opcode_type, 16#0A#),
      2245 => to_slv(opcode_type, 16#0D#),
      2246 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#09#),
      2273 => to_slv(opcode_type, 16#06#),
      2274 => to_slv(opcode_type, 16#02#),
      2275 => to_slv(opcode_type, 16#11#),
      2276 => to_slv(opcode_type, 16#0B#),
      2277 => to_slv(opcode_type, 16#10#),
      2278 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#09#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#03#),
      2307 => to_slv(opcode_type, 16#0B#),
      2308 => to_slv(opcode_type, 16#11#),
      2309 => to_slv(opcode_type, 16#10#),
      2310 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#05#),
      2337 => to_slv(opcode_type, 16#03#),
      2338 => to_slv(opcode_type, 16#07#),
      2339 => to_slv(opcode_type, 16#02#),
      2340 => to_slv(opcode_type, 16#0F#),
      2341 => to_slv(opcode_type, 16#11#),
      2342 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#02#),
      2369 => to_slv(opcode_type, 16#02#),
      2370 => to_slv(opcode_type, 16#07#),
      2371 => to_slv(opcode_type, 16#05#),
      2372 => to_slv(opcode_type, 16#0A#),
      2373 => to_slv(opcode_type, 16#0F#),
      2374 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#05#),
      2401 => to_slv(opcode_type, 16#08#),
      2402 => to_slv(opcode_type, 16#08#),
      2403 => to_slv(opcode_type, 16#0C#),
      2404 => to_slv(opcode_type, 16#0A#),
      2405 => to_slv(opcode_type, 16#0E#),
      2406 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#06#),
      2433 => to_slv(opcode_type, 16#02#),
      2434 => to_slv(opcode_type, 16#06#),
      2435 => to_slv(opcode_type, 16#0D#),
      2436 => to_slv(opcode_type, 16#0A#),
      2437 => to_slv(opcode_type, 16#8E#),
      2438 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#03#),
      2465 => to_slv(opcode_type, 16#04#),
      2466 => to_slv(opcode_type, 16#01#),
      2467 => to_slv(opcode_type, 16#08#),
      2468 => to_slv(opcode_type, 16#10#),
      2469 => to_slv(opcode_type, 16#10#),
      2470 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#04#),
      2497 => to_slv(opcode_type, 16#06#),
      2498 => to_slv(opcode_type, 16#01#),
      2499 => to_slv(opcode_type, 16#05#),
      2500 => to_slv(opcode_type, 16#10#),
      2501 => to_slv(opcode_type, 16#0C#),
      2502 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#02#),
      2529 => to_slv(opcode_type, 16#01#),
      2530 => to_slv(opcode_type, 16#02#),
      2531 => to_slv(opcode_type, 16#08#),
      2532 => to_slv(opcode_type, 16#0C#),
      2533 => to_slv(opcode_type, 16#0C#),
      2534 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#01#),
      2561 => to_slv(opcode_type, 16#08#),
      2562 => to_slv(opcode_type, 16#08#),
      2563 => to_slv(opcode_type, 16#10#),
      2564 => to_slv(opcode_type, 16#0F#),
      2565 => to_slv(opcode_type, 16#0F#),
      2566 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#06#),
      2593 => to_slv(opcode_type, 16#09#),
      2594 => to_slv(opcode_type, 16#03#),
      2595 => to_slv(opcode_type, 16#0E#),
      2596 => to_slv(opcode_type, 16#10#),
      2597 => to_slv(opcode_type, 16#0E#),
      2598 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#04#),
      2625 => to_slv(opcode_type, 16#04#),
      2626 => to_slv(opcode_type, 16#08#),
      2627 => to_slv(opcode_type, 16#02#),
      2628 => to_slv(opcode_type, 16#0C#),
      2629 => to_slv(opcode_type, 16#0B#),
      2630 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#04#),
      2657 => to_slv(opcode_type, 16#05#),
      2658 => to_slv(opcode_type, 16#04#),
      2659 => to_slv(opcode_type, 16#07#),
      2660 => to_slv(opcode_type, 16#10#),
      2661 => to_slv(opcode_type, 16#11#),
      2662 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#03#),
      2689 => to_slv(opcode_type, 16#08#),
      2690 => to_slv(opcode_type, 16#04#),
      2691 => to_slv(opcode_type, 16#05#),
      2692 => to_slv(opcode_type, 16#0A#),
      2693 => to_slv(opcode_type, 16#1A#),
      2694 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#06#),
      2721 => to_slv(opcode_type, 16#06#),
      2722 => to_slv(opcode_type, 16#05#),
      2723 => to_slv(opcode_type, 16#0C#),
      2724 => to_slv(opcode_type, 16#0A#),
      2725 => to_slv(opcode_type, 16#57#),
      2726 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#02#),
      2753 => to_slv(opcode_type, 16#09#),
      2754 => to_slv(opcode_type, 16#03#),
      2755 => to_slv(opcode_type, 16#05#),
      2756 => to_slv(opcode_type, 16#0E#),
      2757 => to_slv(opcode_type, 16#11#),
      2758 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#04#),
      2785 => to_slv(opcode_type, 16#05#),
      2786 => to_slv(opcode_type, 16#03#),
      2787 => to_slv(opcode_type, 16#07#),
      2788 => to_slv(opcode_type, 16#10#),
      2789 => to_slv(opcode_type, 16#0C#),
      2790 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#09#),
      2817 => to_slv(opcode_type, 16#09#),
      2818 => to_slv(opcode_type, 16#01#),
      2819 => to_slv(opcode_type, 16#0E#),
      2820 => to_slv(opcode_type, 16#0E#),
      2821 => to_slv(opcode_type, 16#0F#),
      2822 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#03#),
      2849 => to_slv(opcode_type, 16#06#),
      2850 => to_slv(opcode_type, 16#09#),
      2851 => to_slv(opcode_type, 16#11#),
      2852 => to_slv(opcode_type, 16#37#),
      2853 => to_slv(opcode_type, 16#0D#),
      2854 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#02#),
      2881 => to_slv(opcode_type, 16#09#),
      2882 => to_slv(opcode_type, 16#07#),
      2883 => to_slv(opcode_type, 16#0F#),
      2884 => to_slv(opcode_type, 16#0B#),
      2885 => to_slv(opcode_type, 16#0C#),
      2886 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#04#),
      2913 => to_slv(opcode_type, 16#02#),
      2914 => to_slv(opcode_type, 16#04#),
      2915 => to_slv(opcode_type, 16#06#),
      2916 => to_slv(opcode_type, 16#0A#),
      2917 => to_slv(opcode_type, 16#0A#),
      2918 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#04#),
      2945 => to_slv(opcode_type, 16#08#),
      2946 => to_slv(opcode_type, 16#06#),
      2947 => to_slv(opcode_type, 16#0E#),
      2948 => to_slv(opcode_type, 16#0D#),
      2949 => to_slv(opcode_type, 16#0A#),
      2950 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#04#),
      2977 => to_slv(opcode_type, 16#03#),
      2978 => to_slv(opcode_type, 16#08#),
      2979 => to_slv(opcode_type, 16#04#),
      2980 => to_slv(opcode_type, 16#11#),
      2981 => to_slv(opcode_type, 16#11#),
      2982 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#01#),
      3009 => to_slv(opcode_type, 16#07#),
      3010 => to_slv(opcode_type, 16#08#),
      3011 => to_slv(opcode_type, 16#6D#),
      3012 => to_slv(opcode_type, 16#11#),
      3013 => to_slv(opcode_type, 16#10#),
      3014 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#06#),
      3041 => to_slv(opcode_type, 16#03#),
      3042 => to_slv(opcode_type, 16#06#),
      3043 => to_slv(opcode_type, 16#11#),
      3044 => to_slv(opcode_type, 16#0A#),
      3045 => to_slv(opcode_type, 16#0A#),
      3046 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#01#),
      3073 => to_slv(opcode_type, 16#06#),
      3074 => to_slv(opcode_type, 16#07#),
      3075 => to_slv(opcode_type, 16#0D#),
      3076 => to_slv(opcode_type, 16#11#),
      3077 => to_slv(opcode_type, 16#0B#),
      3078 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#06#),
      3105 => to_slv(opcode_type, 16#03#),
      3106 => to_slv(opcode_type, 16#06#),
      3107 => to_slv(opcode_type, 16#C3#),
      3108 => to_slv(opcode_type, 16#10#),
      3109 => to_slv(opcode_type, 16#41#),
      3110 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#05#),
      3137 => to_slv(opcode_type, 16#09#),
      3138 => to_slv(opcode_type, 16#09#),
      3139 => to_slv(opcode_type, 16#0B#),
      3140 => to_slv(opcode_type, 16#11#),
      3141 => to_slv(opcode_type, 16#0D#),
      3142 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#06#),
      3169 => to_slv(opcode_type, 16#02#),
      3170 => to_slv(opcode_type, 16#06#),
      3171 => to_slv(opcode_type, 16#0A#),
      3172 => to_slv(opcode_type, 16#0F#),
      3173 => to_slv(opcode_type, 16#BA#),
      3174 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#02#),
      3201 => to_slv(opcode_type, 16#01#),
      3202 => to_slv(opcode_type, 16#04#),
      3203 => to_slv(opcode_type, 16#09#),
      3204 => to_slv(opcode_type, 16#11#),
      3205 => to_slv(opcode_type, 16#0D#),
      3206 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#01#),
      3233 => to_slv(opcode_type, 16#04#),
      3234 => to_slv(opcode_type, 16#07#),
      3235 => to_slv(opcode_type, 16#02#),
      3236 => to_slv(opcode_type, 16#11#),
      3237 => to_slv(opcode_type, 16#0D#),
      3238 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#05#),
      3265 => to_slv(opcode_type, 16#01#),
      3266 => to_slv(opcode_type, 16#01#),
      3267 => to_slv(opcode_type, 16#08#),
      3268 => to_slv(opcode_type, 16#1C#),
      3269 => to_slv(opcode_type, 16#0D#),
      3270 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#05#),
      3297 => to_slv(opcode_type, 16#06#),
      3298 => to_slv(opcode_type, 16#05#),
      3299 => to_slv(opcode_type, 16#01#),
      3300 => to_slv(opcode_type, 16#0F#),
      3301 => to_slv(opcode_type, 16#0C#),
      3302 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#01#),
      3329 => to_slv(opcode_type, 16#04#),
      3330 => to_slv(opcode_type, 16#06#),
      3331 => to_slv(opcode_type, 16#05#),
      3332 => to_slv(opcode_type, 16#0B#),
      3333 => to_slv(opcode_type, 16#0B#),
      3334 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#06#),
      3361 => to_slv(opcode_type, 16#06#),
      3362 => to_slv(opcode_type, 16#02#),
      3363 => to_slv(opcode_type, 16#0C#),
      3364 => to_slv(opcode_type, 16#0A#),
      3365 => to_slv(opcode_type, 16#0B#),
      3366 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#07#),
      3393 => to_slv(opcode_type, 16#05#),
      3394 => to_slv(opcode_type, 16#03#),
      3395 => to_slv(opcode_type, 16#04#),
      3396 => to_slv(opcode_type, 16#0B#),
      3397 => to_slv(opcode_type, 16#11#),
      3398 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#06#),
      3425 => to_slv(opcode_type, 16#03#),
      3426 => to_slv(opcode_type, 16#07#),
      3427 => to_slv(opcode_type, 16#0E#),
      3428 => to_slv(opcode_type, 16#53#),
      3429 => to_slv(opcode_type, 16#0A#),
      3430 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#03#),
      3457 => to_slv(opcode_type, 16#01#),
      3458 => to_slv(opcode_type, 16#03#),
      3459 => to_slv(opcode_type, 16#09#),
      3460 => to_slv(opcode_type, 16#0E#),
      3461 => to_slv(opcode_type, 16#11#),
      3462 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#06#),
      3489 => to_slv(opcode_type, 16#07#),
      3490 => to_slv(opcode_type, 16#01#),
      3491 => to_slv(opcode_type, 16#10#),
      3492 => to_slv(opcode_type, 16#0D#),
      3493 => to_slv(opcode_type, 16#0E#),
      3494 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#06#),
      3521 => to_slv(opcode_type, 16#04#),
      3522 => to_slv(opcode_type, 16#04#),
      3523 => to_slv(opcode_type, 16#02#),
      3524 => to_slv(opcode_type, 16#D1#),
      3525 => to_slv(opcode_type, 16#0E#),
      3526 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#07#),
      3553 => to_slv(opcode_type, 16#08#),
      3554 => to_slv(opcode_type, 16#04#),
      3555 => to_slv(opcode_type, 16#0A#),
      3556 => to_slv(opcode_type, 16#11#),
      3557 => to_slv(opcode_type, 16#11#),
      3558 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#01#),
      3585 => to_slv(opcode_type, 16#05#),
      3586 => to_slv(opcode_type, 16#01#),
      3587 => to_slv(opcode_type, 16#06#),
      3588 => to_slv(opcode_type, 16#0D#),
      3589 => to_slv(opcode_type, 16#11#),
      3590 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#05#),
      3617 => to_slv(opcode_type, 16#01#),
      3618 => to_slv(opcode_type, 16#09#),
      3619 => to_slv(opcode_type, 16#02#),
      3620 => to_slv(opcode_type, 16#0E#),
      3621 => to_slv(opcode_type, 16#0E#),
      3622 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#09#),
      3649 => to_slv(opcode_type, 16#09#),
      3650 => to_slv(opcode_type, 16#04#),
      3651 => to_slv(opcode_type, 16#0B#),
      3652 => to_slv(opcode_type, 16#0B#),
      3653 => to_slv(opcode_type, 16#0B#),
      3654 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#03#),
      3681 => to_slv(opcode_type, 16#01#),
      3682 => to_slv(opcode_type, 16#05#),
      3683 => to_slv(opcode_type, 16#07#),
      3684 => to_slv(opcode_type, 16#11#),
      3685 => to_slv(opcode_type, 16#A4#),
      3686 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#08#),
      3713 => to_slv(opcode_type, 16#01#),
      3714 => to_slv(opcode_type, 16#09#),
      3715 => to_slv(opcode_type, 16#11#),
      3716 => to_slv(opcode_type, 16#0F#),
      3717 => to_slv(opcode_type, 16#0E#),
      3718 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#08#),
      3745 => to_slv(opcode_type, 16#02#),
      3746 => to_slv(opcode_type, 16#05#),
      3747 => to_slv(opcode_type, 16#02#),
      3748 => to_slv(opcode_type, 16#0C#),
      3749 => to_slv(opcode_type, 16#0B#),
      3750 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#07#),
      3777 => to_slv(opcode_type, 16#08#),
      3778 => to_slv(opcode_type, 16#05#),
      3779 => to_slv(opcode_type, 16#0D#),
      3780 => to_slv(opcode_type, 16#11#),
      3781 => to_slv(opcode_type, 16#10#),
      3782 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#05#),
      3809 => to_slv(opcode_type, 16#05#),
      3810 => to_slv(opcode_type, 16#01#),
      3811 => to_slv(opcode_type, 16#06#),
      3812 => to_slv(opcode_type, 16#0B#),
      3813 => to_slv(opcode_type, 16#0E#),
      3814 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#02#),
      3841 => to_slv(opcode_type, 16#08#),
      3842 => to_slv(opcode_type, 16#05#),
      3843 => to_slv(opcode_type, 16#01#),
      3844 => to_slv(opcode_type, 16#0C#),
      3845 => to_slv(opcode_type, 16#10#),
      3846 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#08#),
      3873 => to_slv(opcode_type, 16#03#),
      3874 => to_slv(opcode_type, 16#09#),
      3875 => to_slv(opcode_type, 16#0F#),
      3876 => to_slv(opcode_type, 16#0D#),
      3877 => to_slv(opcode_type, 16#0E#),
      3878 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#05#),
      3905 => to_slv(opcode_type, 16#02#),
      3906 => to_slv(opcode_type, 16#03#),
      3907 => to_slv(opcode_type, 16#08#),
      3908 => to_slv(opcode_type, 16#10#),
      3909 => to_slv(opcode_type, 16#0D#),
      3910 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#01#),
      3937 => to_slv(opcode_type, 16#03#),
      3938 => to_slv(opcode_type, 16#09#),
      3939 => to_slv(opcode_type, 16#01#),
      3940 => to_slv(opcode_type, 16#92#),
      3941 => to_slv(opcode_type, 16#10#),
      3942 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#01#),
      3969 => to_slv(opcode_type, 16#09#),
      3970 => to_slv(opcode_type, 16#07#),
      3971 => to_slv(opcode_type, 16#0F#),
      3972 => to_slv(opcode_type, 16#0E#),
      3973 => to_slv(opcode_type, 16#24#),
      3974 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#09#),
      4001 => to_slv(opcode_type, 16#02#),
      4002 => to_slv(opcode_type, 16#03#),
      4003 => to_slv(opcode_type, 16#04#),
      4004 => to_slv(opcode_type, 16#B7#),
      4005 => to_slv(opcode_type, 16#0C#),
      4006 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#09#),
      4033 => to_slv(opcode_type, 16#03#),
      4034 => to_slv(opcode_type, 16#03#),
      4035 => to_slv(opcode_type, 16#02#),
      4036 => to_slv(opcode_type, 16#0D#),
      4037 => to_slv(opcode_type, 16#11#),
      4038 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#05#),
      4065 => to_slv(opcode_type, 16#07#),
      4066 => to_slv(opcode_type, 16#03#),
      4067 => to_slv(opcode_type, 16#02#),
      4068 => to_slv(opcode_type, 16#0F#),
      4069 => to_slv(opcode_type, 16#0E#),
      4070 to 4095 => (others => '0')
  ),

    -- Bin `7`...
    6 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#01#),
      1 => to_slv(opcode_type, 16#04#),
      2 => to_slv(opcode_type, 16#06#),
      3 => to_slv(opcode_type, 16#08#),
      4 => to_slv(opcode_type, 16#6D#),
      5 => to_slv(opcode_type, 16#11#),
      6 => to_slv(opcode_type, 16#0F#),
      7 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#06#),
      33 => to_slv(opcode_type, 16#02#),
      34 => to_slv(opcode_type, 16#07#),
      35 => to_slv(opcode_type, 16#02#),
      36 => to_slv(opcode_type, 16#0A#),
      37 => to_slv(opcode_type, 16#10#),
      38 => to_slv(opcode_type, 16#F7#),
      39 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#04#),
      65 => to_slv(opcode_type, 16#04#),
      66 => to_slv(opcode_type, 16#09#),
      67 => to_slv(opcode_type, 16#02#),
      68 => to_slv(opcode_type, 16#0C#),
      69 => to_slv(opcode_type, 16#02#),
      70 => to_slv(opcode_type, 16#10#),
      71 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#03#),
      97 => to_slv(opcode_type, 16#08#),
      98 => to_slv(opcode_type, 16#07#),
      99 => to_slv(opcode_type, 16#03#),
      100 => to_slv(opcode_type, 16#11#),
      101 => to_slv(opcode_type, 16#0C#),
      102 => to_slv(opcode_type, 16#57#),
      103 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#09#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#03#),
      131 => to_slv(opcode_type, 16#04#),
      132 => to_slv(opcode_type, 16#0A#),
      133 => to_slv(opcode_type, 16#10#),
      134 => to_slv(opcode_type, 16#0A#),
      135 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#01#),
      161 => to_slv(opcode_type, 16#04#),
      162 => to_slv(opcode_type, 16#08#),
      163 => to_slv(opcode_type, 16#04#),
      164 => to_slv(opcode_type, 16#0C#),
      165 => to_slv(opcode_type, 16#04#),
      166 => to_slv(opcode_type, 16#0A#),
      167 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#03#),
      193 => to_slv(opcode_type, 16#02#),
      194 => to_slv(opcode_type, 16#08#),
      195 => to_slv(opcode_type, 16#02#),
      196 => to_slv(opcode_type, 16#11#),
      197 => to_slv(opcode_type, 16#05#),
      198 => to_slv(opcode_type, 16#10#),
      199 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#05#),
      225 => to_slv(opcode_type, 16#05#),
      226 => to_slv(opcode_type, 16#06#),
      227 => to_slv(opcode_type, 16#03#),
      228 => to_slv(opcode_type, 16#0D#),
      229 => to_slv(opcode_type, 16#01#),
      230 => to_slv(opcode_type, 16#12#),
      231 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#09#),
      257 => to_slv(opcode_type, 16#04#),
      258 => to_slv(opcode_type, 16#07#),
      259 => to_slv(opcode_type, 16#03#),
      260 => to_slv(opcode_type, 16#0F#),
      261 => to_slv(opcode_type, 16#68#),
      262 => to_slv(opcode_type, 16#0B#),
      263 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#09#),
      290 => to_slv(opcode_type, 16#03#),
      291 => to_slv(opcode_type, 16#03#),
      292 => to_slv(opcode_type, 16#0B#),
      293 => to_slv(opcode_type, 16#A0#),
      294 => to_slv(opcode_type, 16#0E#),
      295 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#07#),
      321 => to_slv(opcode_type, 16#01#),
      322 => to_slv(opcode_type, 16#09#),
      323 => to_slv(opcode_type, 16#02#),
      324 => to_slv(opcode_type, 16#0F#),
      325 => to_slv(opcode_type, 16#0B#),
      326 => to_slv(opcode_type, 16#0E#),
      327 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#02#),
      353 => to_slv(opcode_type, 16#04#),
      354 => to_slv(opcode_type, 16#06#),
      355 => to_slv(opcode_type, 16#09#),
      356 => to_slv(opcode_type, 16#5F#),
      357 => to_slv(opcode_type, 16#0E#),
      358 => to_slv(opcode_type, 16#0B#),
      359 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#05#),
      385 => to_slv(opcode_type, 16#05#),
      386 => to_slv(opcode_type, 16#06#),
      387 => to_slv(opcode_type, 16#06#),
      388 => to_slv(opcode_type, 16#0F#),
      389 => to_slv(opcode_type, 16#0E#),
      390 => to_slv(opcode_type, 16#0C#),
      391 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#06#),
      417 => to_slv(opcode_type, 16#03#),
      418 => to_slv(opcode_type, 16#05#),
      419 => to_slv(opcode_type, 16#03#),
      420 => to_slv(opcode_type, 16#0B#),
      421 => to_slv(opcode_type, 16#03#),
      422 => to_slv(opcode_type, 16#0C#),
      423 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#08#),
      449 => to_slv(opcode_type, 16#04#),
      450 => to_slv(opcode_type, 16#07#),
      451 => to_slv(opcode_type, 16#01#),
      452 => to_slv(opcode_type, 16#0A#),
      453 => to_slv(opcode_type, 16#0C#),
      454 => to_slv(opcode_type, 16#10#),
      455 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#04#),
      481 => to_slv(opcode_type, 16#02#),
      482 => to_slv(opcode_type, 16#07#),
      483 => to_slv(opcode_type, 16#02#),
      484 => to_slv(opcode_type, 16#0E#),
      485 => to_slv(opcode_type, 16#03#),
      486 => to_slv(opcode_type, 16#11#),
      487 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#08#),
      513 => to_slv(opcode_type, 16#04#),
      514 => to_slv(opcode_type, 16#04#),
      515 => to_slv(opcode_type, 16#05#),
      516 => to_slv(opcode_type, 16#4B#),
      517 => to_slv(opcode_type, 16#01#),
      518 => to_slv(opcode_type, 16#0A#),
      519 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#08#),
      545 => to_slv(opcode_type, 16#01#),
      546 => to_slv(opcode_type, 16#02#),
      547 => to_slv(opcode_type, 16#07#),
      548 => to_slv(opcode_type, 16#0C#),
      549 => to_slv(opcode_type, 16#0C#),
      550 => to_slv(opcode_type, 16#0D#),
      551 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#07#),
      577 => to_slv(opcode_type, 16#02#),
      578 => to_slv(opcode_type, 16#03#),
      579 => to_slv(opcode_type, 16#06#),
      580 => to_slv(opcode_type, 16#0D#),
      581 => to_slv(opcode_type, 16#5D#),
      582 => to_slv(opcode_type, 16#B2#),
      583 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#08#),
      609 => to_slv(opcode_type, 16#05#),
      610 => to_slv(opcode_type, 16#01#),
      611 => to_slv(opcode_type, 16#08#),
      612 => to_slv(opcode_type, 16#0C#),
      613 => to_slv(opcode_type, 16#0B#),
      614 => to_slv(opcode_type, 16#10#),
      615 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#04#),
      641 => to_slv(opcode_type, 16#05#),
      642 => to_slv(opcode_type, 16#07#),
      643 => to_slv(opcode_type, 16#01#),
      644 => to_slv(opcode_type, 16#11#),
      645 => to_slv(opcode_type, 16#04#),
      646 => to_slv(opcode_type, 16#0D#),
      647 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#06#),
      673 => to_slv(opcode_type, 16#03#),
      674 => to_slv(opcode_type, 16#01#),
      675 => to_slv(opcode_type, 16#06#),
      676 => to_slv(opcode_type, 16#0B#),
      677 => to_slv(opcode_type, 16#0A#),
      678 => to_slv(opcode_type, 16#0B#),
      679 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#07#),
      705 => to_slv(opcode_type, 16#04#),
      706 => to_slv(opcode_type, 16#09#),
      707 => to_slv(opcode_type, 16#03#),
      708 => to_slv(opcode_type, 16#0F#),
      709 => to_slv(opcode_type, 16#10#),
      710 => to_slv(opcode_type, 16#0D#),
      711 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#08#),
      737 => to_slv(opcode_type, 16#04#),
      738 => to_slv(opcode_type, 16#09#),
      739 => to_slv(opcode_type, 16#03#),
      740 => to_slv(opcode_type, 16#0E#),
      741 => to_slv(opcode_type, 16#11#),
      742 => to_slv(opcode_type, 16#0E#),
      743 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#06#),
      769 => to_slv(opcode_type, 16#08#),
      770 => to_slv(opcode_type, 16#01#),
      771 => to_slv(opcode_type, 16#04#),
      772 => to_slv(opcode_type, 16#11#),
      773 => to_slv(opcode_type, 16#0E#),
      774 => to_slv(opcode_type, 16#0C#),
      775 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#05#),
      801 => to_slv(opcode_type, 16#09#),
      802 => to_slv(opcode_type, 16#08#),
      803 => to_slv(opcode_type, 16#04#),
      804 => to_slv(opcode_type, 16#10#),
      805 => to_slv(opcode_type, 16#0D#),
      806 => to_slv(opcode_type, 16#0E#),
      807 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#04#),
      833 => to_slv(opcode_type, 16#06#),
      834 => to_slv(opcode_type, 16#06#),
      835 => to_slv(opcode_type, 16#03#),
      836 => to_slv(opcode_type, 16#11#),
      837 => to_slv(opcode_type, 16#11#),
      838 => to_slv(opcode_type, 16#0F#),
      839 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#04#),
      865 => to_slv(opcode_type, 16#09#),
      866 => to_slv(opcode_type, 16#06#),
      867 => to_slv(opcode_type, 16#01#),
      868 => to_slv(opcode_type, 16#C8#),
      869 => to_slv(opcode_type, 16#10#),
      870 => to_slv(opcode_type, 16#0B#),
      871 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#05#),
      897 => to_slv(opcode_type, 16#09#),
      898 => to_slv(opcode_type, 16#01#),
      899 => to_slv(opcode_type, 16#02#),
      900 => to_slv(opcode_type, 16#10#),
      901 => to_slv(opcode_type, 16#03#),
      902 => to_slv(opcode_type, 16#A7#),
      903 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#09#),
      929 => to_slv(opcode_type, 16#01#),
      930 => to_slv(opcode_type, 16#08#),
      931 => to_slv(opcode_type, 16#03#),
      932 => to_slv(opcode_type, 16#0C#),
      933 => to_slv(opcode_type, 16#11#),
      934 => to_slv(opcode_type, 16#10#),
      935 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#04#),
      961 => to_slv(opcode_type, 16#04#),
      962 => to_slv(opcode_type, 16#08#),
      963 => to_slv(opcode_type, 16#05#),
      964 => to_slv(opcode_type, 16#0F#),
      965 => to_slv(opcode_type, 16#05#),
      966 => to_slv(opcode_type, 16#0D#),
      967 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#07#),
      993 => to_slv(opcode_type, 16#09#),
      994 => to_slv(opcode_type, 16#03#),
      995 => to_slv(opcode_type, 16#03#),
      996 => to_slv(opcode_type, 16#11#),
      997 => to_slv(opcode_type, 16#0E#),
      998 => to_slv(opcode_type, 16#AD#),
      999 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#02#),
      1025 => to_slv(opcode_type, 16#04#),
      1026 => to_slv(opcode_type, 16#07#),
      1027 => to_slv(opcode_type, 16#07#),
      1028 => to_slv(opcode_type, 16#0B#),
      1029 => to_slv(opcode_type, 16#10#),
      1030 => to_slv(opcode_type, 16#0C#),
      1031 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#08#),
      1057 => to_slv(opcode_type, 16#07#),
      1058 => to_slv(opcode_type, 16#07#),
      1059 => to_slv(opcode_type, 16#0C#),
      1060 => to_slv(opcode_type, 16#0D#),
      1061 => to_slv(opcode_type, 16#0E#),
      1062 => to_slv(opcode_type, 16#10#),
      1063 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#01#),
      1089 => to_slv(opcode_type, 16#06#),
      1090 => to_slv(opcode_type, 16#09#),
      1091 => to_slv(opcode_type, 16#03#),
      1092 => to_slv(opcode_type, 16#0B#),
      1093 => to_slv(opcode_type, 16#F0#),
      1094 => to_slv(opcode_type, 16#0D#),
      1095 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#05#),
      1121 => to_slv(opcode_type, 16#05#),
      1122 => to_slv(opcode_type, 16#07#),
      1123 => to_slv(opcode_type, 16#04#),
      1124 => to_slv(opcode_type, 16#63#),
      1125 => to_slv(opcode_type, 16#02#),
      1126 => to_slv(opcode_type, 16#0D#),
      1127 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#01#),
      1153 => to_slv(opcode_type, 16#06#),
      1154 => to_slv(opcode_type, 16#09#),
      1155 => to_slv(opcode_type, 16#02#),
      1156 => to_slv(opcode_type, 16#0F#),
      1157 => to_slv(opcode_type, 16#0D#),
      1158 => to_slv(opcode_type, 16#0F#),
      1159 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#03#),
      1185 => to_slv(opcode_type, 16#05#),
      1186 => to_slv(opcode_type, 16#07#),
      1187 => to_slv(opcode_type, 16#09#),
      1188 => to_slv(opcode_type, 16#0E#),
      1189 => to_slv(opcode_type, 16#0A#),
      1190 => to_slv(opcode_type, 16#0E#),
      1191 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#07#),
      1217 => to_slv(opcode_type, 16#03#),
      1218 => to_slv(opcode_type, 16#01#),
      1219 => to_slv(opcode_type, 16#03#),
      1220 => to_slv(opcode_type, 16#0B#),
      1221 => to_slv(opcode_type, 16#02#),
      1222 => to_slv(opcode_type, 16#0F#),
      1223 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#07#),
      1249 => to_slv(opcode_type, 16#07#),
      1250 => to_slv(opcode_type, 16#04#),
      1251 => to_slv(opcode_type, 16#01#),
      1252 => to_slv(opcode_type, 16#0F#),
      1253 => to_slv(opcode_type, 16#0C#),
      1254 => to_slv(opcode_type, 16#0E#),
      1255 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#05#),
      1281 => to_slv(opcode_type, 16#01#),
      1282 => to_slv(opcode_type, 16#08#),
      1283 => to_slv(opcode_type, 16#05#),
      1284 => to_slv(opcode_type, 16#0C#),
      1285 => to_slv(opcode_type, 16#03#),
      1286 => to_slv(opcode_type, 16#0D#),
      1287 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#01#),
      1313 => to_slv(opcode_type, 16#06#),
      1314 => to_slv(opcode_type, 16#06#),
      1315 => to_slv(opcode_type, 16#02#),
      1316 => to_slv(opcode_type, 16#6E#),
      1317 => to_slv(opcode_type, 16#0A#),
      1318 => to_slv(opcode_type, 16#5C#),
      1319 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#02#),
      1345 => to_slv(opcode_type, 16#05#),
      1346 => to_slv(opcode_type, 16#08#),
      1347 => to_slv(opcode_type, 16#06#),
      1348 => to_slv(opcode_type, 16#2D#),
      1349 => to_slv(opcode_type, 16#0E#),
      1350 => to_slv(opcode_type, 16#51#),
      1351 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#06#),
      1377 => to_slv(opcode_type, 16#02#),
      1378 => to_slv(opcode_type, 16#02#),
      1379 => to_slv(opcode_type, 16#07#),
      1380 => to_slv(opcode_type, 16#0F#),
      1381 => to_slv(opcode_type, 16#10#),
      1382 => to_slv(opcode_type, 16#0D#),
      1383 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#07#),
      1409 => to_slv(opcode_type, 16#08#),
      1410 => to_slv(opcode_type, 16#05#),
      1411 => to_slv(opcode_type, 16#05#),
      1412 => to_slv(opcode_type, 16#0C#),
      1413 => to_slv(opcode_type, 16#0A#),
      1414 => to_slv(opcode_type, 16#0A#),
      1415 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#06#),
      1441 => to_slv(opcode_type, 16#07#),
      1442 => to_slv(opcode_type, 16#07#),
      1443 => to_slv(opcode_type, 16#0B#),
      1444 => to_slv(opcode_type, 16#0B#),
      1445 => to_slv(opcode_type, 16#0D#),
      1446 => to_slv(opcode_type, 16#0D#),
      1447 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#04#),
      1473 => to_slv(opcode_type, 16#02#),
      1474 => to_slv(opcode_type, 16#07#),
      1475 => to_slv(opcode_type, 16#05#),
      1476 => to_slv(opcode_type, 16#0C#),
      1477 => to_slv(opcode_type, 16#03#),
      1478 => to_slv(opcode_type, 16#0C#),
      1479 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#03#),
      1505 => to_slv(opcode_type, 16#02#),
      1506 => to_slv(opcode_type, 16#06#),
      1507 => to_slv(opcode_type, 16#05#),
      1508 => to_slv(opcode_type, 16#0B#),
      1509 => to_slv(opcode_type, 16#04#),
      1510 => to_slv(opcode_type, 16#0B#),
      1511 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#04#),
      1537 => to_slv(opcode_type, 16#03#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#02#),
      1540 => to_slv(opcode_type, 16#0C#),
      1541 => to_slv(opcode_type, 16#02#),
      1542 => to_slv(opcode_type, 16#0F#),
      1543 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#02#),
      1569 => to_slv(opcode_type, 16#05#),
      1570 => to_slv(opcode_type, 16#07#),
      1571 => to_slv(opcode_type, 16#05#),
      1572 => to_slv(opcode_type, 16#0A#),
      1573 => to_slv(opcode_type, 16#02#),
      1574 => to_slv(opcode_type, 16#0E#),
      1575 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#07#),
      1601 => to_slv(opcode_type, 16#09#),
      1602 => to_slv(opcode_type, 16#02#),
      1603 => to_slv(opcode_type, 16#04#),
      1604 => to_slv(opcode_type, 16#0A#),
      1605 => to_slv(opcode_type, 16#19#),
      1606 => to_slv(opcode_type, 16#0B#),
      1607 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#04#),
      1633 => to_slv(opcode_type, 16#06#),
      1634 => to_slv(opcode_type, 16#06#),
      1635 => to_slv(opcode_type, 16#04#),
      1636 => to_slv(opcode_type, 16#0D#),
      1637 => to_slv(opcode_type, 16#0B#),
      1638 => to_slv(opcode_type, 16#0C#),
      1639 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#06#),
      1665 => to_slv(opcode_type, 16#02#),
      1666 => to_slv(opcode_type, 16#03#),
      1667 => to_slv(opcode_type, 16#08#),
      1668 => to_slv(opcode_type, 16#0F#),
      1669 => to_slv(opcode_type, 16#10#),
      1670 => to_slv(opcode_type, 16#97#),
      1671 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#03#),
      1697 => to_slv(opcode_type, 16#01#),
      1698 => to_slv(opcode_type, 16#08#),
      1699 => to_slv(opcode_type, 16#08#),
      1700 => to_slv(opcode_type, 16#0B#),
      1701 => to_slv(opcode_type, 16#0D#),
      1702 => to_slv(opcode_type, 16#9A#),
      1703 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#05#),
      1729 => to_slv(opcode_type, 16#05#),
      1730 => to_slv(opcode_type, 16#08#),
      1731 => to_slv(opcode_type, 16#06#),
      1732 => to_slv(opcode_type, 16#0D#),
      1733 => to_slv(opcode_type, 16#0A#),
      1734 => to_slv(opcode_type, 16#89#),
      1735 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#02#),
      1761 => to_slv(opcode_type, 16#07#),
      1762 => to_slv(opcode_type, 16#09#),
      1763 => to_slv(opcode_type, 16#01#),
      1764 => to_slv(opcode_type, 16#11#),
      1765 => to_slv(opcode_type, 16#11#),
      1766 => to_slv(opcode_type, 16#0E#),
      1767 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#06#),
      1793 => to_slv(opcode_type, 16#09#),
      1794 => to_slv(opcode_type, 16#07#),
      1795 => to_slv(opcode_type, 16#10#),
      1796 => to_slv(opcode_type, 16#10#),
      1797 => to_slv(opcode_type, 16#0B#),
      1798 => to_slv(opcode_type, 16#A9#),
      1799 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#05#),
      1825 => to_slv(opcode_type, 16#06#),
      1826 => to_slv(opcode_type, 16#05#),
      1827 => to_slv(opcode_type, 16#09#),
      1828 => to_slv(opcode_type, 16#0E#),
      1829 => to_slv(opcode_type, 16#12#),
      1830 => to_slv(opcode_type, 16#10#),
      1831 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#06#),
      1857 => to_slv(opcode_type, 16#05#),
      1858 => to_slv(opcode_type, 16#07#),
      1859 => to_slv(opcode_type, 16#05#),
      1860 => to_slv(opcode_type, 16#0C#),
      1861 => to_slv(opcode_type, 16#0F#),
      1862 => to_slv(opcode_type, 16#AB#),
      1863 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#09#),
      1889 => to_slv(opcode_type, 16#09#),
      1890 => to_slv(opcode_type, 16#03#),
      1891 => to_slv(opcode_type, 16#04#),
      1892 => to_slv(opcode_type, 16#11#),
      1893 => to_slv(opcode_type, 16#95#),
      1894 => to_slv(opcode_type, 16#11#),
      1895 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#06#),
      1921 => to_slv(opcode_type, 16#07#),
      1922 => to_slv(opcode_type, 16#01#),
      1923 => to_slv(opcode_type, 16#02#),
      1924 => to_slv(opcode_type, 16#0F#),
      1925 => to_slv(opcode_type, 16#0B#),
      1926 => to_slv(opcode_type, 16#0A#),
      1927 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#04#),
      1953 => to_slv(opcode_type, 16#05#),
      1954 => to_slv(opcode_type, 16#08#),
      1955 => to_slv(opcode_type, 16#07#),
      1956 => to_slv(opcode_type, 16#0D#),
      1957 => to_slv(opcode_type, 16#11#),
      1958 => to_slv(opcode_type, 16#0B#),
      1959 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#08#),
      1985 => to_slv(opcode_type, 16#03#),
      1986 => to_slv(opcode_type, 16#04#),
      1987 => to_slv(opcode_type, 16#09#),
      1988 => to_slv(opcode_type, 16#0D#),
      1989 => to_slv(opcode_type, 16#11#),
      1990 => to_slv(opcode_type, 16#0F#),
      1991 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#07#),
      2017 => to_slv(opcode_type, 16#04#),
      2018 => to_slv(opcode_type, 16#02#),
      2019 => to_slv(opcode_type, 16#07#),
      2020 => to_slv(opcode_type, 16#10#),
      2021 => to_slv(opcode_type, 16#11#),
      2022 => to_slv(opcode_type, 16#0A#),
      2023 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#07#),
      2049 => to_slv(opcode_type, 16#03#),
      2050 => to_slv(opcode_type, 16#05#),
      2051 => to_slv(opcode_type, 16#06#),
      2052 => to_slv(opcode_type, 16#11#),
      2053 => to_slv(opcode_type, 16#0F#),
      2054 => to_slv(opcode_type, 16#0B#),
      2055 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#08#),
      2081 => to_slv(opcode_type, 16#03#),
      2082 => to_slv(opcode_type, 16#07#),
      2083 => to_slv(opcode_type, 16#04#),
      2084 => to_slv(opcode_type, 16#0D#),
      2085 => to_slv(opcode_type, 16#10#),
      2086 => to_slv(opcode_type, 16#26#),
      2087 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#05#),
      2113 => to_slv(opcode_type, 16#05#),
      2114 => to_slv(opcode_type, 16#06#),
      2115 => to_slv(opcode_type, 16#07#),
      2116 => to_slv(opcode_type, 16#0F#),
      2117 => to_slv(opcode_type, 16#0E#),
      2118 => to_slv(opcode_type, 16#10#),
      2119 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#02#),
      2145 => to_slv(opcode_type, 16#02#),
      2146 => to_slv(opcode_type, 16#07#),
      2147 => to_slv(opcode_type, 16#05#),
      2148 => to_slv(opcode_type, 16#0E#),
      2149 => to_slv(opcode_type, 16#04#),
      2150 => to_slv(opcode_type, 16#11#),
      2151 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#04#),
      2177 => to_slv(opcode_type, 16#07#),
      2178 => to_slv(opcode_type, 16#08#),
      2179 => to_slv(opcode_type, 16#03#),
      2180 => to_slv(opcode_type, 16#0C#),
      2181 => to_slv(opcode_type, 16#0F#),
      2182 => to_slv(opcode_type, 16#11#),
      2183 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#03#),
      2209 => to_slv(opcode_type, 16#07#),
      2210 => to_slv(opcode_type, 16#03#),
      2211 => to_slv(opcode_type, 16#09#),
      2212 => to_slv(opcode_type, 16#0B#),
      2213 => to_slv(opcode_type, 16#11#),
      2214 => to_slv(opcode_type, 16#11#),
      2215 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#05#),
      2241 => to_slv(opcode_type, 16#03#),
      2242 => to_slv(opcode_type, 16#08#),
      2243 => to_slv(opcode_type, 16#06#),
      2244 => to_slv(opcode_type, 16#0D#),
      2245 => to_slv(opcode_type, 16#0B#),
      2246 => to_slv(opcode_type, 16#0B#),
      2247 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#03#),
      2273 => to_slv(opcode_type, 16#05#),
      2274 => to_slv(opcode_type, 16#08#),
      2275 => to_slv(opcode_type, 16#09#),
      2276 => to_slv(opcode_type, 16#0F#),
      2277 => to_slv(opcode_type, 16#10#),
      2278 => to_slv(opcode_type, 16#0F#),
      2279 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#02#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#09#),
      2307 => to_slv(opcode_type, 16#01#),
      2308 => to_slv(opcode_type, 16#0F#),
      2309 => to_slv(opcode_type, 16#0D#),
      2310 => to_slv(opcode_type, 16#0D#),
      2311 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#08#),
      2337 => to_slv(opcode_type, 16#01#),
      2338 => to_slv(opcode_type, 16#07#),
      2339 => to_slv(opcode_type, 16#05#),
      2340 => to_slv(opcode_type, 16#0C#),
      2341 => to_slv(opcode_type, 16#99#),
      2342 => to_slv(opcode_type, 16#10#),
      2343 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#04#),
      2369 => to_slv(opcode_type, 16#03#),
      2370 => to_slv(opcode_type, 16#07#),
      2371 => to_slv(opcode_type, 16#07#),
      2372 => to_slv(opcode_type, 16#10#),
      2373 => to_slv(opcode_type, 16#0E#),
      2374 => to_slv(opcode_type, 16#0D#),
      2375 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#08#),
      2401 => to_slv(opcode_type, 16#04#),
      2402 => to_slv(opcode_type, 16#07#),
      2403 => to_slv(opcode_type, 16#04#),
      2404 => to_slv(opcode_type, 16#0F#),
      2405 => to_slv(opcode_type, 16#0A#),
      2406 => to_slv(opcode_type, 16#0A#),
      2407 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#02#),
      2433 => to_slv(opcode_type, 16#05#),
      2434 => to_slv(opcode_type, 16#09#),
      2435 => to_slv(opcode_type, 16#07#),
      2436 => to_slv(opcode_type, 16#0C#),
      2437 => to_slv(opcode_type, 16#0C#),
      2438 => to_slv(opcode_type, 16#0E#),
      2439 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#05#),
      2465 => to_slv(opcode_type, 16#08#),
      2466 => to_slv(opcode_type, 16#08#),
      2467 => to_slv(opcode_type, 16#03#),
      2468 => to_slv(opcode_type, 16#81#),
      2469 => to_slv(opcode_type, 16#11#),
      2470 => to_slv(opcode_type, 16#10#),
      2471 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#06#),
      2497 => to_slv(opcode_type, 16#02#),
      2498 => to_slv(opcode_type, 16#08#),
      2499 => to_slv(opcode_type, 16#02#),
      2500 => to_slv(opcode_type, 16#10#),
      2501 => to_slv(opcode_type, 16#0C#),
      2502 => to_slv(opcode_type, 16#10#),
      2503 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#01#),
      2529 => to_slv(opcode_type, 16#08#),
      2530 => to_slv(opcode_type, 16#09#),
      2531 => to_slv(opcode_type, 16#03#),
      2532 => to_slv(opcode_type, 16#0C#),
      2533 => to_slv(opcode_type, 16#0A#),
      2534 => to_slv(opcode_type, 16#0B#),
      2535 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#04#),
      2561 => to_slv(opcode_type, 16#08#),
      2562 => to_slv(opcode_type, 16#04#),
      2563 => to_slv(opcode_type, 16#01#),
      2564 => to_slv(opcode_type, 16#11#),
      2565 => to_slv(opcode_type, 16#03#),
      2566 => to_slv(opcode_type, 16#0E#),
      2567 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#03#),
      2593 => to_slv(opcode_type, 16#03#),
      2594 => to_slv(opcode_type, 16#06#),
      2595 => to_slv(opcode_type, 16#08#),
      2596 => to_slv(opcode_type, 16#11#),
      2597 => to_slv(opcode_type, 16#0E#),
      2598 => to_slv(opcode_type, 16#11#),
      2599 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#07#),
      2625 => to_slv(opcode_type, 16#09#),
      2626 => to_slv(opcode_type, 16#04#),
      2627 => to_slv(opcode_type, 16#01#),
      2628 => to_slv(opcode_type, 16#0B#),
      2629 => to_slv(opcode_type, 16#0A#),
      2630 => to_slv(opcode_type, 16#3A#),
      2631 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#09#),
      2657 => to_slv(opcode_type, 16#03#),
      2658 => to_slv(opcode_type, 16#09#),
      2659 => to_slv(opcode_type, 16#03#),
      2660 => to_slv(opcode_type, 16#0E#),
      2661 => to_slv(opcode_type, 16#11#),
      2662 => to_slv(opcode_type, 16#0C#),
      2663 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#04#),
      2689 => to_slv(opcode_type, 16#09#),
      2690 => to_slv(opcode_type, 16#03#),
      2691 => to_slv(opcode_type, 16#07#),
      2692 => to_slv(opcode_type, 16#11#),
      2693 => to_slv(opcode_type, 16#0F#),
      2694 => to_slv(opcode_type, 16#11#),
      2695 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#06#),
      2721 => to_slv(opcode_type, 16#04#),
      2722 => to_slv(opcode_type, 16#09#),
      2723 => to_slv(opcode_type, 16#01#),
      2724 => to_slv(opcode_type, 16#0F#),
      2725 => to_slv(opcode_type, 16#0E#),
      2726 => to_slv(opcode_type, 16#0F#),
      2727 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#04#),
      2753 => to_slv(opcode_type, 16#09#),
      2754 => to_slv(opcode_type, 16#01#),
      2755 => to_slv(opcode_type, 16#04#),
      2756 => to_slv(opcode_type, 16#10#),
      2757 => to_slv(opcode_type, 16#04#),
      2758 => to_slv(opcode_type, 16#0E#),
      2759 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#02#),
      2785 => to_slv(opcode_type, 16#06#),
      2786 => to_slv(opcode_type, 16#02#),
      2787 => to_slv(opcode_type, 16#02#),
      2788 => to_slv(opcode_type, 16#0E#),
      2789 => to_slv(opcode_type, 16#03#),
      2790 => to_slv(opcode_type, 16#AC#),
      2791 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#02#),
      2817 => to_slv(opcode_type, 16#05#),
      2818 => to_slv(opcode_type, 16#08#),
      2819 => to_slv(opcode_type, 16#05#),
      2820 => to_slv(opcode_type, 16#11#),
      2821 => to_slv(opcode_type, 16#02#),
      2822 => to_slv(opcode_type, 16#0B#),
      2823 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#05#),
      2849 => to_slv(opcode_type, 16#05#),
      2850 => to_slv(opcode_type, 16#08#),
      2851 => to_slv(opcode_type, 16#01#),
      2852 => to_slv(opcode_type, 16#0B#),
      2853 => to_slv(opcode_type, 16#02#),
      2854 => to_slv(opcode_type, 16#10#),
      2855 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#03#),
      2881 => to_slv(opcode_type, 16#05#),
      2882 => to_slv(opcode_type, 16#07#),
      2883 => to_slv(opcode_type, 16#01#),
      2884 => to_slv(opcode_type, 16#11#),
      2885 => to_slv(opcode_type, 16#01#),
      2886 => to_slv(opcode_type, 16#0A#),
      2887 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#04#),
      2913 => to_slv(opcode_type, 16#04#),
      2914 => to_slv(opcode_type, 16#09#),
      2915 => to_slv(opcode_type, 16#08#),
      2916 => to_slv(opcode_type, 16#0E#),
      2917 => to_slv(opcode_type, 16#87#),
      2918 => to_slv(opcode_type, 16#0C#),
      2919 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#04#),
      2945 => to_slv(opcode_type, 16#05#),
      2946 => to_slv(opcode_type, 16#08#),
      2947 => to_slv(opcode_type, 16#01#),
      2948 => to_slv(opcode_type, 16#0D#),
      2949 => to_slv(opcode_type, 16#02#),
      2950 => to_slv(opcode_type, 16#28#),
      2951 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#04#),
      2977 => to_slv(opcode_type, 16#03#),
      2978 => to_slv(opcode_type, 16#07#),
      2979 => to_slv(opcode_type, 16#08#),
      2980 => to_slv(opcode_type, 16#0D#),
      2981 => to_slv(opcode_type, 16#0E#),
      2982 => to_slv(opcode_type, 16#0B#),
      2983 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#05#),
      3009 => to_slv(opcode_type, 16#01#),
      3010 => to_slv(opcode_type, 16#09#),
      3011 => to_slv(opcode_type, 16#05#),
      3012 => to_slv(opcode_type, 16#0F#),
      3013 => to_slv(opcode_type, 16#02#),
      3014 => to_slv(opcode_type, 16#0D#),
      3015 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#01#),
      3041 => to_slv(opcode_type, 16#04#),
      3042 => to_slv(opcode_type, 16#08#),
      3043 => to_slv(opcode_type, 16#03#),
      3044 => to_slv(opcode_type, 16#0B#),
      3045 => to_slv(opcode_type, 16#05#),
      3046 => to_slv(opcode_type, 16#0C#),
      3047 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#07#),
      3073 => to_slv(opcode_type, 16#07#),
      3074 => to_slv(opcode_type, 16#03#),
      3075 => to_slv(opcode_type, 16#03#),
      3076 => to_slv(opcode_type, 16#0C#),
      3077 => to_slv(opcode_type, 16#10#),
      3078 => to_slv(opcode_type, 16#61#),
      3079 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#02#),
      3105 => to_slv(opcode_type, 16#02#),
      3106 => to_slv(opcode_type, 16#09#),
      3107 => to_slv(opcode_type, 16#09#),
      3108 => to_slv(opcode_type, 16#10#),
      3109 => to_slv(opcode_type, 16#0E#),
      3110 => to_slv(opcode_type, 16#0B#),
      3111 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#02#),
      3137 => to_slv(opcode_type, 16#06#),
      3138 => to_slv(opcode_type, 16#01#),
      3139 => to_slv(opcode_type, 16#03#),
      3140 => to_slv(opcode_type, 16#0B#),
      3141 => to_slv(opcode_type, 16#04#),
      3142 => to_slv(opcode_type, 16#10#),
      3143 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#05#),
      3169 => to_slv(opcode_type, 16#06#),
      3170 => to_slv(opcode_type, 16#01#),
      3171 => to_slv(opcode_type, 16#05#),
      3172 => to_slv(opcode_type, 16#EB#),
      3173 => to_slv(opcode_type, 16#02#),
      3174 => to_slv(opcode_type, 16#0B#),
      3175 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#05#),
      3201 => to_slv(opcode_type, 16#04#),
      3202 => to_slv(opcode_type, 16#08#),
      3203 => to_slv(opcode_type, 16#03#),
      3204 => to_slv(opcode_type, 16#0C#),
      3205 => to_slv(opcode_type, 16#01#),
      3206 => to_slv(opcode_type, 16#0E#),
      3207 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#04#),
      3234 => to_slv(opcode_type, 16#06#),
      3235 => to_slv(opcode_type, 16#01#),
      3236 => to_slv(opcode_type, 16#0D#),
      3237 => to_slv(opcode_type, 16#0A#),
      3238 => to_slv(opcode_type, 16#0F#),
      3239 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#01#),
      3265 => to_slv(opcode_type, 16#01#),
      3266 => to_slv(opcode_type, 16#08#),
      3267 => to_slv(opcode_type, 16#01#),
      3268 => to_slv(opcode_type, 16#10#),
      3269 => to_slv(opcode_type, 16#01#),
      3270 => to_slv(opcode_type, 16#10#),
      3271 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#07#),
      3297 => to_slv(opcode_type, 16#07#),
      3298 => to_slv(opcode_type, 16#08#),
      3299 => to_slv(opcode_type, 16#11#),
      3300 => to_slv(opcode_type, 16#0E#),
      3301 => to_slv(opcode_type, 16#49#),
      3302 => to_slv(opcode_type, 16#10#),
      3303 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#06#),
      3329 => to_slv(opcode_type, 16#08#),
      3330 => to_slv(opcode_type, 16#09#),
      3331 => to_slv(opcode_type, 16#0F#),
      3332 => to_slv(opcode_type, 16#0B#),
      3333 => to_slv(opcode_type, 16#11#),
      3334 => to_slv(opcode_type, 16#0C#),
      3335 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#05#),
      3361 => to_slv(opcode_type, 16#07#),
      3362 => to_slv(opcode_type, 16#06#),
      3363 => to_slv(opcode_type, 16#01#),
      3364 => to_slv(opcode_type, 16#0E#),
      3365 => to_slv(opcode_type, 16#11#),
      3366 => to_slv(opcode_type, 16#10#),
      3367 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#08#),
      3393 => to_slv(opcode_type, 16#01#),
      3394 => to_slv(opcode_type, 16#01#),
      3395 => to_slv(opcode_type, 16#02#),
      3396 => to_slv(opcode_type, 16#0A#),
      3397 => to_slv(opcode_type, 16#01#),
      3398 => to_slv(opcode_type, 16#3E#),
      3399 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#07#),
      3426 => to_slv(opcode_type, 16#09#),
      3427 => to_slv(opcode_type, 16#0A#),
      3428 => to_slv(opcode_type, 16#0C#),
      3429 => to_slv(opcode_type, 16#11#),
      3430 => to_slv(opcode_type, 16#0C#),
      3431 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#04#),
      3457 => to_slv(opcode_type, 16#07#),
      3458 => to_slv(opcode_type, 16#09#),
      3459 => to_slv(opcode_type, 16#02#),
      3460 => to_slv(opcode_type, 16#0C#),
      3461 => to_slv(opcode_type, 16#0D#),
      3462 => to_slv(opcode_type, 16#0B#),
      3463 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#07#),
      3489 => to_slv(opcode_type, 16#05#),
      3490 => to_slv(opcode_type, 16#06#),
      3491 => to_slv(opcode_type, 16#01#),
      3492 => to_slv(opcode_type, 16#0E#),
      3493 => to_slv(opcode_type, 16#0C#),
      3494 => to_slv(opcode_type, 16#48#),
      3495 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#06#),
      3521 => to_slv(opcode_type, 16#09#),
      3522 => to_slv(opcode_type, 16#02#),
      3523 => to_slv(opcode_type, 16#05#),
      3524 => to_slv(opcode_type, 16#0E#),
      3525 => to_slv(opcode_type, 16#0C#),
      3526 => to_slv(opcode_type, 16#10#),
      3527 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#06#),
      3553 => to_slv(opcode_type, 16#06#),
      3554 => to_slv(opcode_type, 16#04#),
      3555 => to_slv(opcode_type, 16#04#),
      3556 => to_slv(opcode_type, 16#0F#),
      3557 => to_slv(opcode_type, 16#18#),
      3558 => to_slv(opcode_type, 16#0E#),
      3559 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#05#),
      3585 => to_slv(opcode_type, 16#07#),
      3586 => to_slv(opcode_type, 16#05#),
      3587 => to_slv(opcode_type, 16#07#),
      3588 => to_slv(opcode_type, 16#0D#),
      3589 => to_slv(opcode_type, 16#10#),
      3590 => to_slv(opcode_type, 16#0B#),
      3591 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#01#),
      3617 => to_slv(opcode_type, 16#05#),
      3618 => to_slv(opcode_type, 16#06#),
      3619 => to_slv(opcode_type, 16#08#),
      3620 => to_slv(opcode_type, 16#0E#),
      3621 => to_slv(opcode_type, 16#0D#),
      3622 => to_slv(opcode_type, 16#0F#),
      3623 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#05#),
      3649 => to_slv(opcode_type, 16#07#),
      3650 => to_slv(opcode_type, 16#07#),
      3651 => to_slv(opcode_type, 16#05#),
      3652 => to_slv(opcode_type, 16#10#),
      3653 => to_slv(opcode_type, 16#0B#),
      3654 => to_slv(opcode_type, 16#0A#),
      3655 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#03#),
      3681 => to_slv(opcode_type, 16#05#),
      3682 => to_slv(opcode_type, 16#09#),
      3683 => to_slv(opcode_type, 16#09#),
      3684 => to_slv(opcode_type, 16#0F#),
      3685 => to_slv(opcode_type, 16#11#),
      3686 => to_slv(opcode_type, 16#0D#),
      3687 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#04#),
      3713 => to_slv(opcode_type, 16#05#),
      3714 => to_slv(opcode_type, 16#07#),
      3715 => to_slv(opcode_type, 16#04#),
      3716 => to_slv(opcode_type, 16#0C#),
      3717 => to_slv(opcode_type, 16#01#),
      3718 => to_slv(opcode_type, 16#10#),
      3719 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#02#),
      3745 => to_slv(opcode_type, 16#04#),
      3746 => to_slv(opcode_type, 16#09#),
      3747 => to_slv(opcode_type, 16#03#),
      3748 => to_slv(opcode_type, 16#10#),
      3749 => to_slv(opcode_type, 16#04#),
      3750 => to_slv(opcode_type, 16#50#),
      3751 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#03#),
      3777 => to_slv(opcode_type, 16#04#),
      3778 => to_slv(opcode_type, 16#07#),
      3779 => to_slv(opcode_type, 16#07#),
      3780 => to_slv(opcode_type, 16#0A#),
      3781 => to_slv(opcode_type, 16#0E#),
      3782 => to_slv(opcode_type, 16#0C#),
      3783 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#09#),
      3809 => to_slv(opcode_type, 16#06#),
      3810 => to_slv(opcode_type, 16#02#),
      3811 => to_slv(opcode_type, 16#02#),
      3812 => to_slv(opcode_type, 16#0D#),
      3813 => to_slv(opcode_type, 16#0E#),
      3814 => to_slv(opcode_type, 16#0B#),
      3815 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#04#),
      3841 => to_slv(opcode_type, 16#04#),
      3842 => to_slv(opcode_type, 16#09#),
      3843 => to_slv(opcode_type, 16#04#),
      3844 => to_slv(opcode_type, 16#0D#),
      3845 => to_slv(opcode_type, 16#03#),
      3846 => to_slv(opcode_type, 16#10#),
      3847 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#06#),
      3873 => to_slv(opcode_type, 16#07#),
      3874 => to_slv(opcode_type, 16#08#),
      3875 => to_slv(opcode_type, 16#0B#),
      3876 => to_slv(opcode_type, 16#11#),
      3877 => to_slv(opcode_type, 16#0D#),
      3878 => to_slv(opcode_type, 16#6C#),
      3879 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#05#),
      3905 => to_slv(opcode_type, 16#09#),
      3906 => to_slv(opcode_type, 16#07#),
      3907 => to_slv(opcode_type, 16#03#),
      3908 => to_slv(opcode_type, 16#0C#),
      3909 => to_slv(opcode_type, 16#0F#),
      3910 => to_slv(opcode_type, 16#0A#),
      3911 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#05#),
      3937 => to_slv(opcode_type, 16#01#),
      3938 => to_slv(opcode_type, 16#06#),
      3939 => to_slv(opcode_type, 16#08#),
      3940 => to_slv(opcode_type, 16#12#),
      3941 => to_slv(opcode_type, 16#0B#),
      3942 => to_slv(opcode_type, 16#11#),
      3943 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#03#),
      3969 => to_slv(opcode_type, 16#08#),
      3970 => to_slv(opcode_type, 16#05#),
      3971 => to_slv(opcode_type, 16#05#),
      3972 => to_slv(opcode_type, 16#0F#),
      3973 => to_slv(opcode_type, 16#02#),
      3974 => to_slv(opcode_type, 16#11#),
      3975 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#01#),
      4001 => to_slv(opcode_type, 16#03#),
      4002 => to_slv(opcode_type, 16#07#),
      4003 => to_slv(opcode_type, 16#07#),
      4004 => to_slv(opcode_type, 16#0E#),
      4005 => to_slv(opcode_type, 16#0C#),
      4006 => to_slv(opcode_type, 16#0A#),
      4007 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#04#),
      4033 => to_slv(opcode_type, 16#08#),
      4034 => to_slv(opcode_type, 16#02#),
      4035 => to_slv(opcode_type, 16#06#),
      4036 => to_slv(opcode_type, 16#0D#),
      4037 => to_slv(opcode_type, 16#11#),
      4038 => to_slv(opcode_type, 16#2F#),
      4039 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#01#),
      4065 => to_slv(opcode_type, 16#03#),
      4066 => to_slv(opcode_type, 16#08#),
      4067 => to_slv(opcode_type, 16#07#),
      4068 => to_slv(opcode_type, 16#0B#),
      4069 => to_slv(opcode_type, 16#0B#),
      4070 => to_slv(opcode_type, 16#0D#),
      4071 to 4095 => (others => '0')
  ),

    -- Bin `8`...
    7 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#06#),
      1 => to_slv(opcode_type, 16#08#),
      2 => to_slv(opcode_type, 16#02#),
      3 => to_slv(opcode_type, 16#01#),
      4 => to_slv(opcode_type, 16#0F#),
      5 => to_slv(opcode_type, 16#03#),
      6 => to_slv(opcode_type, 16#0E#),
      7 => to_slv(opcode_type, 16#11#),
      8 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#07#),
      33 => to_slv(opcode_type, 16#06#),
      34 => to_slv(opcode_type, 16#03#),
      35 => to_slv(opcode_type, 16#03#),
      36 => to_slv(opcode_type, 16#0F#),
      37 => to_slv(opcode_type, 16#04#),
      38 => to_slv(opcode_type, 16#0E#),
      39 => to_slv(opcode_type, 16#10#),
      40 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#02#),
      65 => to_slv(opcode_type, 16#01#),
      66 => to_slv(opcode_type, 16#09#),
      67 => to_slv(opcode_type, 16#04#),
      68 => to_slv(opcode_type, 16#10#),
      69 => to_slv(opcode_type, 16#08#),
      70 => to_slv(opcode_type, 16#11#),
      71 => to_slv(opcode_type, 16#0E#),
      72 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#02#),
      97 => to_slv(opcode_type, 16#06#),
      98 => to_slv(opcode_type, 16#07#),
      99 => to_slv(opcode_type, 16#07#),
      100 => to_slv(opcode_type, 16#11#),
      101 => to_slv(opcode_type, 16#0A#),
      102 => to_slv(opcode_type, 16#0D#),
      103 => to_slv(opcode_type, 16#0E#),
      104 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#04#),
      129 => to_slv(opcode_type, 16#06#),
      130 => to_slv(opcode_type, 16#08#),
      131 => to_slv(opcode_type, 16#01#),
      132 => to_slv(opcode_type, 16#0A#),
      133 => to_slv(opcode_type, 16#05#),
      134 => to_slv(opcode_type, 16#11#),
      135 => to_slv(opcode_type, 16#C3#),
      136 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#09#),
      161 => to_slv(opcode_type, 16#07#),
      162 => to_slv(opcode_type, 16#07#),
      163 => to_slv(opcode_type, 16#04#),
      164 => to_slv(opcode_type, 16#0E#),
      165 => to_slv(opcode_type, 16#0E#),
      166 => to_slv(opcode_type, 16#0E#),
      167 => to_slv(opcode_type, 16#10#),
      168 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#09#),
      193 => to_slv(opcode_type, 16#08#),
      194 => to_slv(opcode_type, 16#03#),
      195 => to_slv(opcode_type, 16#01#),
      196 => to_slv(opcode_type, 16#0E#),
      197 => to_slv(opcode_type, 16#01#),
      198 => to_slv(opcode_type, 16#90#),
      199 => to_slv(opcode_type, 16#10#),
      200 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#04#),
      225 => to_slv(opcode_type, 16#06#),
      226 => to_slv(opcode_type, 16#01#),
      227 => to_slv(opcode_type, 16#03#),
      228 => to_slv(opcode_type, 16#0D#),
      229 => to_slv(opcode_type, 16#05#),
      230 => to_slv(opcode_type, 16#02#),
      231 => to_slv(opcode_type, 16#0E#),
      232 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#05#),
      257 => to_slv(opcode_type, 16#01#),
      258 => to_slv(opcode_type, 16#07#),
      259 => to_slv(opcode_type, 16#08#),
      260 => to_slv(opcode_type, 16#0B#),
      261 => to_slv(opcode_type, 16#14#),
      262 => to_slv(opcode_type, 16#04#),
      263 => to_slv(opcode_type, 16#0B#),
      264 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#03#),
      290 => to_slv(opcode_type, 16#03#),
      291 => to_slv(opcode_type, 16#01#),
      292 => to_slv(opcode_type, 16#0E#),
      293 => to_slv(opcode_type, 16#01#),
      294 => to_slv(opcode_type, 16#01#),
      295 => to_slv(opcode_type, 16#0F#),
      296 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#03#),
      321 => to_slv(opcode_type, 16#09#),
      322 => to_slv(opcode_type, 16#03#),
      323 => to_slv(opcode_type, 16#01#),
      324 => to_slv(opcode_type, 16#0E#),
      325 => to_slv(opcode_type, 16#08#),
      326 => to_slv(opcode_type, 16#24#),
      327 => to_slv(opcode_type, 16#0D#),
      328 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#09#),
      353 => to_slv(opcode_type, 16#07#),
      354 => to_slv(opcode_type, 16#03#),
      355 => to_slv(opcode_type, 16#09#),
      356 => to_slv(opcode_type, 16#11#),
      357 => to_slv(opcode_type, 16#B9#),
      358 => to_slv(opcode_type, 16#0B#),
      359 => to_slv(opcode_type, 16#0C#),
      360 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#01#),
      385 => to_slv(opcode_type, 16#05#),
      386 => to_slv(opcode_type, 16#06#),
      387 => to_slv(opcode_type, 16#04#),
      388 => to_slv(opcode_type, 16#0F#),
      389 => to_slv(opcode_type, 16#09#),
      390 => to_slv(opcode_type, 16#0D#),
      391 => to_slv(opcode_type, 16#0F#),
      392 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#08#),
      417 => to_slv(opcode_type, 16#08#),
      418 => to_slv(opcode_type, 16#01#),
      419 => to_slv(opcode_type, 16#05#),
      420 => to_slv(opcode_type, 16#0D#),
      421 => to_slv(opcode_type, 16#05#),
      422 => to_slv(opcode_type, 16#0A#),
      423 => to_slv(opcode_type, 16#0F#),
      424 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#07#),
      449 => to_slv(opcode_type, 16#08#),
      450 => to_slv(opcode_type, 16#03#),
      451 => to_slv(opcode_type, 16#01#),
      452 => to_slv(opcode_type, 16#0B#),
      453 => to_slv(opcode_type, 16#03#),
      454 => to_slv(opcode_type, 16#0A#),
      455 => to_slv(opcode_type, 16#0E#),
      456 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#01#),
      481 => to_slv(opcode_type, 16#02#),
      482 => to_slv(opcode_type, 16#09#),
      483 => to_slv(opcode_type, 16#08#),
      484 => to_slv(opcode_type, 16#D1#),
      485 => to_slv(opcode_type, 16#0F#),
      486 => to_slv(opcode_type, 16#01#),
      487 => to_slv(opcode_type, 16#0E#),
      488 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#05#),
      513 => to_slv(opcode_type, 16#04#),
      514 => to_slv(opcode_type, 16#07#),
      515 => to_slv(opcode_type, 16#06#),
      516 => to_slv(opcode_type, 16#0C#),
      517 => to_slv(opcode_type, 16#11#),
      518 => to_slv(opcode_type, 16#04#),
      519 => to_slv(opcode_type, 16#0E#),
      520 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#02#),
      545 => to_slv(opcode_type, 16#05#),
      546 => to_slv(opcode_type, 16#08#),
      547 => to_slv(opcode_type, 16#09#),
      548 => to_slv(opcode_type, 16#0F#),
      549 => to_slv(opcode_type, 16#0C#),
      550 => to_slv(opcode_type, 16#02#),
      551 => to_slv(opcode_type, 16#0A#),
      552 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#09#),
      577 => to_slv(opcode_type, 16#05#),
      578 => to_slv(opcode_type, 16#06#),
      579 => to_slv(opcode_type, 16#03#),
      580 => to_slv(opcode_type, 16#0C#),
      581 => to_slv(opcode_type, 16#02#),
      582 => to_slv(opcode_type, 16#8E#),
      583 => to_slv(opcode_type, 16#0F#),
      584 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#09#),
      609 => to_slv(opcode_type, 16#03#),
      610 => to_slv(opcode_type, 16#07#),
      611 => to_slv(opcode_type, 16#02#),
      612 => to_slv(opcode_type, 16#0B#),
      613 => to_slv(opcode_type, 16#03#),
      614 => to_slv(opcode_type, 16#0A#),
      615 => to_slv(opcode_type, 16#0A#),
      616 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#01#),
      641 => to_slv(opcode_type, 16#03#),
      642 => to_slv(opcode_type, 16#06#),
      643 => to_slv(opcode_type, 16#08#),
      644 => to_slv(opcode_type, 16#0B#),
      645 => to_slv(opcode_type, 16#11#),
      646 => to_slv(opcode_type, 16#02#),
      647 => to_slv(opcode_type, 16#0B#),
      648 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#03#),
      673 => to_slv(opcode_type, 16#08#),
      674 => to_slv(opcode_type, 16#02#),
      675 => to_slv(opcode_type, 16#09#),
      676 => to_slv(opcode_type, 16#0C#),
      677 => to_slv(opcode_type, 16#0A#),
      678 => to_slv(opcode_type, 16#05#),
      679 => to_slv(opcode_type, 16#10#),
      680 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#08#),
      705 => to_slv(opcode_type, 16#04#),
      706 => to_slv(opcode_type, 16#01#),
      707 => to_slv(opcode_type, 16#03#),
      708 => to_slv(opcode_type, 16#0E#),
      709 => to_slv(opcode_type, 16#03#),
      710 => to_slv(opcode_type, 16#01#),
      711 => to_slv(opcode_type, 16#41#),
      712 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#06#),
      737 => to_slv(opcode_type, 16#03#),
      738 => to_slv(opcode_type, 16#08#),
      739 => to_slv(opcode_type, 16#05#),
      740 => to_slv(opcode_type, 16#0A#),
      741 => to_slv(opcode_type, 16#05#),
      742 => to_slv(opcode_type, 16#0B#),
      743 => to_slv(opcode_type, 16#0E#),
      744 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#02#),
      769 => to_slv(opcode_type, 16#07#),
      770 => to_slv(opcode_type, 16#06#),
      771 => to_slv(opcode_type, 16#02#),
      772 => to_slv(opcode_type, 16#10#),
      773 => to_slv(opcode_type, 16#04#),
      774 => to_slv(opcode_type, 16#11#),
      775 => to_slv(opcode_type, 16#FB#),
      776 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#06#),
      801 => to_slv(opcode_type, 16#04#),
      802 => to_slv(opcode_type, 16#02#),
      803 => to_slv(opcode_type, 16#07#),
      804 => to_slv(opcode_type, 16#0F#),
      805 => to_slv(opcode_type, 16#0A#),
      806 => to_slv(opcode_type, 16#03#),
      807 => to_slv(opcode_type, 16#0A#),
      808 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#03#),
      833 => to_slv(opcode_type, 16#09#),
      834 => to_slv(opcode_type, 16#03#),
      835 => to_slv(opcode_type, 16#07#),
      836 => to_slv(opcode_type, 16#0F#),
      837 => to_slv(opcode_type, 16#0E#),
      838 => to_slv(opcode_type, 16#04#),
      839 => to_slv(opcode_type, 16#0C#),
      840 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#09#),
      865 => to_slv(opcode_type, 16#08#),
      866 => to_slv(opcode_type, 16#05#),
      867 => to_slv(opcode_type, 16#09#),
      868 => to_slv(opcode_type, 16#53#),
      869 => to_slv(opcode_type, 16#0B#),
      870 => to_slv(opcode_type, 16#0E#),
      871 => to_slv(opcode_type, 16#0D#),
      872 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#06#),
      897 => to_slv(opcode_type, 16#09#),
      898 => to_slv(opcode_type, 16#01#),
      899 => to_slv(opcode_type, 16#08#),
      900 => to_slv(opcode_type, 16#0C#),
      901 => to_slv(opcode_type, 16#D2#),
      902 => to_slv(opcode_type, 16#0C#),
      903 => to_slv(opcode_type, 16#0A#),
      904 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#02#),
      929 => to_slv(opcode_type, 16#02#),
      930 => to_slv(opcode_type, 16#07#),
      931 => to_slv(opcode_type, 16#01#),
      932 => to_slv(opcode_type, 16#0E#),
      933 => to_slv(opcode_type, 16#06#),
      934 => to_slv(opcode_type, 16#10#),
      935 => to_slv(opcode_type, 16#0D#),
      936 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#05#),
      961 => to_slv(opcode_type, 16#02#),
      962 => to_slv(opcode_type, 16#07#),
      963 => to_slv(opcode_type, 16#08#),
      964 => to_slv(opcode_type, 16#10#),
      965 => to_slv(opcode_type, 16#0E#),
      966 => to_slv(opcode_type, 16#02#),
      967 => to_slv(opcode_type, 16#11#),
      968 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#05#),
      993 => to_slv(opcode_type, 16#02#),
      994 => to_slv(opcode_type, 16#06#),
      995 => to_slv(opcode_type, 16#07#),
      996 => to_slv(opcode_type, 16#10#),
      997 => to_slv(opcode_type, 16#0E#),
      998 => to_slv(opcode_type, 16#04#),
      999 => to_slv(opcode_type, 16#76#),
      1000 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#05#),
      1025 => to_slv(opcode_type, 16#06#),
      1026 => to_slv(opcode_type, 16#02#),
      1027 => to_slv(opcode_type, 16#07#),
      1028 => to_slv(opcode_type, 16#0B#),
      1029 => to_slv(opcode_type, 16#0A#),
      1030 => to_slv(opcode_type, 16#02#),
      1031 => to_slv(opcode_type, 16#11#),
      1032 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#01#),
      1057 => to_slv(opcode_type, 16#09#),
      1058 => to_slv(opcode_type, 16#02#),
      1059 => to_slv(opcode_type, 16#08#),
      1060 => to_slv(opcode_type, 16#0E#),
      1061 => to_slv(opcode_type, 16#11#),
      1062 => to_slv(opcode_type, 16#05#),
      1063 => to_slv(opcode_type, 16#0A#),
      1064 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#08#),
      1089 => to_slv(opcode_type, 16#04#),
      1090 => to_slv(opcode_type, 16#06#),
      1091 => to_slv(opcode_type, 16#05#),
      1092 => to_slv(opcode_type, 16#0F#),
      1093 => to_slv(opcode_type, 16#02#),
      1094 => to_slv(opcode_type, 16#0A#),
      1095 => to_slv(opcode_type, 16#0E#),
      1096 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#06#),
      1121 => to_slv(opcode_type, 16#03#),
      1122 => to_slv(opcode_type, 16#05#),
      1123 => to_slv(opcode_type, 16#04#),
      1124 => to_slv(opcode_type, 16#0E#),
      1125 => to_slv(opcode_type, 16#03#),
      1126 => to_slv(opcode_type, 16#02#),
      1127 => to_slv(opcode_type, 16#0F#),
      1128 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#09#),
      1153 => to_slv(opcode_type, 16#09#),
      1154 => to_slv(opcode_type, 16#07#),
      1155 => to_slv(opcode_type, 16#01#),
      1156 => to_slv(opcode_type, 16#0D#),
      1157 => to_slv(opcode_type, 16#0E#),
      1158 => to_slv(opcode_type, 16#0C#),
      1159 => to_slv(opcode_type, 16#0F#),
      1160 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#01#),
      1185 => to_slv(opcode_type, 16#08#),
      1186 => to_slv(opcode_type, 16#01#),
      1187 => to_slv(opcode_type, 16#03#),
      1188 => to_slv(opcode_type, 16#0F#),
      1189 => to_slv(opcode_type, 16#01#),
      1190 => to_slv(opcode_type, 16#03#),
      1191 => to_slv(opcode_type, 16#0B#),
      1192 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#05#),
      1217 => to_slv(opcode_type, 16#07#),
      1218 => to_slv(opcode_type, 16#08#),
      1219 => to_slv(opcode_type, 16#09#),
      1220 => to_slv(opcode_type, 16#0A#),
      1221 => to_slv(opcode_type, 16#74#),
      1222 => to_slv(opcode_type, 16#0B#),
      1223 => to_slv(opcode_type, 16#0F#),
      1224 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#08#),
      1249 => to_slv(opcode_type, 16#09#),
      1250 => to_slv(opcode_type, 16#08#),
      1251 => to_slv(opcode_type, 16#02#),
      1252 => to_slv(opcode_type, 16#10#),
      1253 => to_slv(opcode_type, 16#0E#),
      1254 => to_slv(opcode_type, 16#0A#),
      1255 => to_slv(opcode_type, 16#11#),
      1256 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#03#),
      1281 => to_slv(opcode_type, 16#05#),
      1282 => to_slv(opcode_type, 16#07#),
      1283 => to_slv(opcode_type, 16#06#),
      1284 => to_slv(opcode_type, 16#0C#),
      1285 => to_slv(opcode_type, 16#10#),
      1286 => to_slv(opcode_type, 16#01#),
      1287 => to_slv(opcode_type, 16#11#),
      1288 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#01#),
      1313 => to_slv(opcode_type, 16#08#),
      1314 => to_slv(opcode_type, 16#08#),
      1315 => to_slv(opcode_type, 16#05#),
      1316 => to_slv(opcode_type, 16#0C#),
      1317 => to_slv(opcode_type, 16#02#),
      1318 => to_slv(opcode_type, 16#0C#),
      1319 => to_slv(opcode_type, 16#0F#),
      1320 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#01#),
      1345 => to_slv(opcode_type, 16#01#),
      1346 => to_slv(opcode_type, 16#09#),
      1347 => to_slv(opcode_type, 16#09#),
      1348 => to_slv(opcode_type, 16#0C#),
      1349 => to_slv(opcode_type, 16#0B#),
      1350 => to_slv(opcode_type, 16#04#),
      1351 => to_slv(opcode_type, 16#F7#),
      1352 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#07#),
      1377 => to_slv(opcode_type, 16#01#),
      1378 => to_slv(opcode_type, 16#06#),
      1379 => to_slv(opcode_type, 16#07#),
      1380 => to_slv(opcode_type, 16#0E#),
      1381 => to_slv(opcode_type, 16#8B#),
      1382 => to_slv(opcode_type, 16#33#),
      1383 => to_slv(opcode_type, 16#0F#),
      1384 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#02#),
      1409 => to_slv(opcode_type, 16#02#),
      1410 => to_slv(opcode_type, 16#07#),
      1411 => to_slv(opcode_type, 16#08#),
      1412 => to_slv(opcode_type, 16#11#),
      1413 => to_slv(opcode_type, 16#0D#),
      1414 => to_slv(opcode_type, 16#02#),
      1415 => to_slv(opcode_type, 16#0F#),
      1416 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#02#),
      1441 => to_slv(opcode_type, 16#08#),
      1442 => to_slv(opcode_type, 16#08#),
      1443 => to_slv(opcode_type, 16#07#),
      1444 => to_slv(opcode_type, 16#11#),
      1445 => to_slv(opcode_type, 16#0D#),
      1446 => to_slv(opcode_type, 16#0E#),
      1447 => to_slv(opcode_type, 16#0C#),
      1448 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#03#),
      1473 => to_slv(opcode_type, 16#01#),
      1474 => to_slv(opcode_type, 16#06#),
      1475 => to_slv(opcode_type, 16#08#),
      1476 => to_slv(opcode_type, 16#0E#),
      1477 => to_slv(opcode_type, 16#0B#),
      1478 => to_slv(opcode_type, 16#04#),
      1479 => to_slv(opcode_type, 16#11#),
      1480 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#06#),
      1505 => to_slv(opcode_type, 16#02#),
      1506 => to_slv(opcode_type, 16#08#),
      1507 => to_slv(opcode_type, 16#03#),
      1508 => to_slv(opcode_type, 16#0E#),
      1509 => to_slv(opcode_type, 16#03#),
      1510 => to_slv(opcode_type, 16#0E#),
      1511 => to_slv(opcode_type, 16#10#),
      1512 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#05#),
      1537 => to_slv(opcode_type, 16#07#),
      1538 => to_slv(opcode_type, 16#02#),
      1539 => to_slv(opcode_type, 16#05#),
      1540 => to_slv(opcode_type, 16#0F#),
      1541 => to_slv(opcode_type, 16#01#),
      1542 => to_slv(opcode_type, 16#04#),
      1543 => to_slv(opcode_type, 16#0E#),
      1544 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#02#),
      1569 => to_slv(opcode_type, 16#02#),
      1570 => to_slv(opcode_type, 16#07#),
      1571 => to_slv(opcode_type, 16#05#),
      1572 => to_slv(opcode_type, 16#0C#),
      1573 => to_slv(opcode_type, 16#06#),
      1574 => to_slv(opcode_type, 16#FD#),
      1575 => to_slv(opcode_type, 16#0F#),
      1576 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#02#),
      1601 => to_slv(opcode_type, 16#03#),
      1602 => to_slv(opcode_type, 16#07#),
      1603 => to_slv(opcode_type, 16#08#),
      1604 => to_slv(opcode_type, 16#0B#),
      1605 => to_slv(opcode_type, 16#D5#),
      1606 => to_slv(opcode_type, 16#04#),
      1607 => to_slv(opcode_type, 16#0C#),
      1608 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#01#),
      1633 => to_slv(opcode_type, 16#08#),
      1634 => to_slv(opcode_type, 16#06#),
      1635 => to_slv(opcode_type, 16#04#),
      1636 => to_slv(opcode_type, 16#11#),
      1637 => to_slv(opcode_type, 16#01#),
      1638 => to_slv(opcode_type, 16#11#),
      1639 => to_slv(opcode_type, 16#0A#),
      1640 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#04#),
      1666 => to_slv(opcode_type, 16#08#),
      1667 => to_slv(opcode_type, 16#02#),
      1668 => to_slv(opcode_type, 16#0A#),
      1669 => to_slv(opcode_type, 16#05#),
      1670 => to_slv(opcode_type, 16#0A#),
      1671 => to_slv(opcode_type, 16#0C#),
      1672 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#04#),
      1697 => to_slv(opcode_type, 16#01#),
      1698 => to_slv(opcode_type, 16#09#),
      1699 => to_slv(opcode_type, 16#08#),
      1700 => to_slv(opcode_type, 16#D5#),
      1701 => to_slv(opcode_type, 16#0A#),
      1702 => to_slv(opcode_type, 16#02#),
      1703 => to_slv(opcode_type, 16#0C#),
      1704 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#03#),
      1729 => to_slv(opcode_type, 16#05#),
      1730 => to_slv(opcode_type, 16#07#),
      1731 => to_slv(opcode_type, 16#08#),
      1732 => to_slv(opcode_type, 16#10#),
      1733 => to_slv(opcode_type, 16#0A#),
      1734 => to_slv(opcode_type, 16#01#),
      1735 => to_slv(opcode_type, 16#0C#),
      1736 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#01#),
      1761 => to_slv(opcode_type, 16#03#),
      1762 => to_slv(opcode_type, 16#07#),
      1763 => to_slv(opcode_type, 16#07#),
      1764 => to_slv(opcode_type, 16#11#),
      1765 => to_slv(opcode_type, 16#10#),
      1766 => to_slv(opcode_type, 16#03#),
      1767 => to_slv(opcode_type, 16#10#),
      1768 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#03#),
      1793 => to_slv(opcode_type, 16#01#),
      1794 => to_slv(opcode_type, 16#07#),
      1795 => to_slv(opcode_type, 16#04#),
      1796 => to_slv(opcode_type, 16#0B#),
      1797 => to_slv(opcode_type, 16#07#),
      1798 => to_slv(opcode_type, 16#10#),
      1799 => to_slv(opcode_type, 16#0A#),
      1800 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#05#),
      1825 => to_slv(opcode_type, 16#02#),
      1826 => to_slv(opcode_type, 16#06#),
      1827 => to_slv(opcode_type, 16#08#),
      1828 => to_slv(opcode_type, 16#0A#),
      1829 => to_slv(opcode_type, 16#0F#),
      1830 => to_slv(opcode_type, 16#03#),
      1831 => to_slv(opcode_type, 16#0B#),
      1832 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#09#),
      1857 => to_slv(opcode_type, 16#04#),
      1858 => to_slv(opcode_type, 16#05#),
      1859 => to_slv(opcode_type, 16#07#),
      1860 => to_slv(opcode_type, 16#11#),
      1861 => to_slv(opcode_type, 16#B9#),
      1862 => to_slv(opcode_type, 16#02#),
      1863 => to_slv(opcode_type, 16#0C#),
      1864 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#08#),
      1889 => to_slv(opcode_type, 16#08#),
      1890 => to_slv(opcode_type, 16#08#),
      1891 => to_slv(opcode_type, 16#01#),
      1892 => to_slv(opcode_type, 16#10#),
      1893 => to_slv(opcode_type, 16#0C#),
      1894 => to_slv(opcode_type, 16#0A#),
      1895 => to_slv(opcode_type, 16#0A#),
      1896 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#08#),
      1921 => to_slv(opcode_type, 16#05#),
      1922 => to_slv(opcode_type, 16#05#),
      1923 => to_slv(opcode_type, 16#07#),
      1924 => to_slv(opcode_type, 16#49#),
      1925 => to_slv(opcode_type, 16#0A#),
      1926 => to_slv(opcode_type, 16#01#),
      1927 => to_slv(opcode_type, 16#0C#),
      1928 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#03#),
      1953 => to_slv(opcode_type, 16#07#),
      1954 => to_slv(opcode_type, 16#05#),
      1955 => to_slv(opcode_type, 16#02#),
      1956 => to_slv(opcode_type, 16#0E#),
      1957 => to_slv(opcode_type, 16#09#),
      1958 => to_slv(opcode_type, 16#0A#),
      1959 => to_slv(opcode_type, 16#0B#),
      1960 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#08#),
      1985 => to_slv(opcode_type, 16#07#),
      1986 => to_slv(opcode_type, 16#01#),
      1987 => to_slv(opcode_type, 16#03#),
      1988 => to_slv(opcode_type, 16#0C#),
      1989 => to_slv(opcode_type, 16#01#),
      1990 => to_slv(opcode_type, 16#0B#),
      1991 => to_slv(opcode_type, 16#0D#),
      1992 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#08#),
      2017 => to_slv(opcode_type, 16#02#),
      2018 => to_slv(opcode_type, 16#05#),
      2019 => to_slv(opcode_type, 16#01#),
      2020 => to_slv(opcode_type, 16#0B#),
      2021 => to_slv(opcode_type, 16#04#),
      2022 => to_slv(opcode_type, 16#02#),
      2023 => to_slv(opcode_type, 16#0D#),
      2024 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#01#),
      2049 => to_slv(opcode_type, 16#05#),
      2050 => to_slv(opcode_type, 16#08#),
      2051 => to_slv(opcode_type, 16#08#),
      2052 => to_slv(opcode_type, 16#AC#),
      2053 => to_slv(opcode_type, 16#0F#),
      2054 => to_slv(opcode_type, 16#02#),
      2055 => to_slv(opcode_type, 16#10#),
      2056 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#09#),
      2081 => to_slv(opcode_type, 16#07#),
      2082 => to_slv(opcode_type, 16#07#),
      2083 => to_slv(opcode_type, 16#05#),
      2084 => to_slv(opcode_type, 16#11#),
      2085 => to_slv(opcode_type, 16#11#),
      2086 => to_slv(opcode_type, 16#10#),
      2087 => to_slv(opcode_type, 16#28#),
      2088 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#01#),
      2113 => to_slv(opcode_type, 16#07#),
      2114 => to_slv(opcode_type, 16#08#),
      2115 => to_slv(opcode_type, 16#08#),
      2116 => to_slv(opcode_type, 16#0A#),
      2117 => to_slv(opcode_type, 16#11#),
      2118 => to_slv(opcode_type, 16#0D#),
      2119 => to_slv(opcode_type, 16#11#),
      2120 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#07#),
      2146 => to_slv(opcode_type, 16#05#),
      2147 => to_slv(opcode_type, 16#08#),
      2148 => to_slv(opcode_type, 16#0C#),
      2149 => to_slv(opcode_type, 16#0D#),
      2150 => to_slv(opcode_type, 16#11#),
      2151 => to_slv(opcode_type, 16#0F#),
      2152 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#03#),
      2177 => to_slv(opcode_type, 16#04#),
      2178 => to_slv(opcode_type, 16#07#),
      2179 => to_slv(opcode_type, 16#06#),
      2180 => to_slv(opcode_type, 16#0E#),
      2181 => to_slv(opcode_type, 16#0B#),
      2182 => to_slv(opcode_type, 16#02#),
      2183 => to_slv(opcode_type, 16#0F#),
      2184 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#01#),
      2209 => to_slv(opcode_type, 16#02#),
      2210 => to_slv(opcode_type, 16#09#),
      2211 => to_slv(opcode_type, 16#09#),
      2212 => to_slv(opcode_type, 16#0B#),
      2213 => to_slv(opcode_type, 16#0B#),
      2214 => to_slv(opcode_type, 16#04#),
      2215 => to_slv(opcode_type, 16#0C#),
      2216 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#07#),
      2241 => to_slv(opcode_type, 16#06#),
      2242 => to_slv(opcode_type, 16#07#),
      2243 => to_slv(opcode_type, 16#05#),
      2244 => to_slv(opcode_type, 16#0D#),
      2245 => to_slv(opcode_type, 16#0B#),
      2246 => to_slv(opcode_type, 16#0E#),
      2247 => to_slv(opcode_type, 16#0B#),
      2248 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#09#),
      2273 => to_slv(opcode_type, 16#08#),
      2274 => to_slv(opcode_type, 16#04#),
      2275 => to_slv(opcode_type, 16#02#),
      2276 => to_slv(opcode_type, 16#0B#),
      2277 => to_slv(opcode_type, 16#05#),
      2278 => to_slv(opcode_type, 16#0D#),
      2279 => to_slv(opcode_type, 16#0C#),
      2280 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#05#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#09#),
      2307 => to_slv(opcode_type, 16#08#),
      2308 => to_slv(opcode_type, 16#0D#),
      2309 => to_slv(opcode_type, 16#0C#),
      2310 => to_slv(opcode_type, 16#0C#),
      2311 => to_slv(opcode_type, 16#11#),
      2312 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#05#),
      2337 => to_slv(opcode_type, 16#08#),
      2338 => to_slv(opcode_type, 16#07#),
      2339 => to_slv(opcode_type, 16#03#),
      2340 => to_slv(opcode_type, 16#10#),
      2341 => to_slv(opcode_type, 16#01#),
      2342 => to_slv(opcode_type, 16#0A#),
      2343 => to_slv(opcode_type, 16#0F#),
      2344 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#08#),
      2369 => to_slv(opcode_type, 16#06#),
      2370 => to_slv(opcode_type, 16#09#),
      2371 => to_slv(opcode_type, 16#01#),
      2372 => to_slv(opcode_type, 16#84#),
      2373 => to_slv(opcode_type, 16#10#),
      2374 => to_slv(opcode_type, 16#11#),
      2375 => to_slv(opcode_type, 16#10#),
      2376 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#04#),
      2401 => to_slv(opcode_type, 16#04#),
      2402 => to_slv(opcode_type, 16#08#),
      2403 => to_slv(opcode_type, 16#05#),
      2404 => to_slv(opcode_type, 16#0F#),
      2405 => to_slv(opcode_type, 16#09#),
      2406 => to_slv(opcode_type, 16#0B#),
      2407 => to_slv(opcode_type, 16#0E#),
      2408 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#02#),
      2433 => to_slv(opcode_type, 16#08#),
      2434 => to_slv(opcode_type, 16#01#),
      2435 => to_slv(opcode_type, 16#08#),
      2436 => to_slv(opcode_type, 16#0C#),
      2437 => to_slv(opcode_type, 16#0C#),
      2438 => to_slv(opcode_type, 16#02#),
      2439 => to_slv(opcode_type, 16#0E#),
      2440 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#03#),
      2465 => to_slv(opcode_type, 16#08#),
      2466 => to_slv(opcode_type, 16#08#),
      2467 => to_slv(opcode_type, 16#02#),
      2468 => to_slv(opcode_type, 16#0B#),
      2469 => to_slv(opcode_type, 16#01#),
      2470 => to_slv(opcode_type, 16#0E#),
      2471 => to_slv(opcode_type, 16#0D#),
      2472 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#01#),
      2497 => to_slv(opcode_type, 16#04#),
      2498 => to_slv(opcode_type, 16#09#),
      2499 => to_slv(opcode_type, 16#09#),
      2500 => to_slv(opcode_type, 16#10#),
      2501 => to_slv(opcode_type, 16#0A#),
      2502 => to_slv(opcode_type, 16#05#),
      2503 => to_slv(opcode_type, 16#AF#),
      2504 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#03#),
      2529 => to_slv(opcode_type, 16#04#),
      2530 => to_slv(opcode_type, 16#08#),
      2531 => to_slv(opcode_type, 16#06#),
      2532 => to_slv(opcode_type, 16#0C#),
      2533 => to_slv(opcode_type, 16#0B#),
      2534 => to_slv(opcode_type, 16#02#),
      2535 => to_slv(opcode_type, 16#0C#),
      2536 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#08#),
      2561 => to_slv(opcode_type, 16#01#),
      2562 => to_slv(opcode_type, 16#08#),
      2563 => to_slv(opcode_type, 16#05#),
      2564 => to_slv(opcode_type, 16#79#),
      2565 => to_slv(opcode_type, 16#04#),
      2566 => to_slv(opcode_type, 16#0C#),
      2567 => to_slv(opcode_type, 16#0D#),
      2568 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#05#),
      2593 => to_slv(opcode_type, 16#01#),
      2594 => to_slv(opcode_type, 16#06#),
      2595 => to_slv(opcode_type, 16#05#),
      2596 => to_slv(opcode_type, 16#0D#),
      2597 => to_slv(opcode_type, 16#07#),
      2598 => to_slv(opcode_type, 16#0F#),
      2599 => to_slv(opcode_type, 16#0E#),
      2600 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#09#),
      2625 => to_slv(opcode_type, 16#06#),
      2626 => to_slv(opcode_type, 16#06#),
      2627 => to_slv(opcode_type, 16#01#),
      2628 => to_slv(opcode_type, 16#42#),
      2629 => to_slv(opcode_type, 16#0D#),
      2630 => to_slv(opcode_type, 16#5B#),
      2631 => to_slv(opcode_type, 16#0E#),
      2632 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#03#),
      2657 => to_slv(opcode_type, 16#02#),
      2658 => to_slv(opcode_type, 16#06#),
      2659 => to_slv(opcode_type, 16#08#),
      2660 => to_slv(opcode_type, 16#0E#),
      2661 => to_slv(opcode_type, 16#0D#),
      2662 => to_slv(opcode_type, 16#01#),
      2663 => to_slv(opcode_type, 16#0B#),
      2664 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#06#),
      2689 => to_slv(opcode_type, 16#09#),
      2690 => to_slv(opcode_type, 16#06#),
      2691 => to_slv(opcode_type, 16#03#),
      2692 => to_slv(opcode_type, 16#0A#),
      2693 => to_slv(opcode_type, 16#0E#),
      2694 => to_slv(opcode_type, 16#4F#),
      2695 => to_slv(opcode_type, 16#0B#),
      2696 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#05#),
      2721 => to_slv(opcode_type, 16#06#),
      2722 => to_slv(opcode_type, 16#02#),
      2723 => to_slv(opcode_type, 16#05#),
      2724 => to_slv(opcode_type, 16#0E#),
      2725 => to_slv(opcode_type, 16#05#),
      2726 => to_slv(opcode_type, 16#03#),
      2727 => to_slv(opcode_type, 16#9A#),
      2728 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#09#),
      2753 => to_slv(opcode_type, 16#09#),
      2754 => to_slv(opcode_type, 16#06#),
      2755 => to_slv(opcode_type, 16#03#),
      2756 => to_slv(opcode_type, 16#0C#),
      2757 => to_slv(opcode_type, 16#0A#),
      2758 => to_slv(opcode_type, 16#11#),
      2759 => to_slv(opcode_type, 16#0C#),
      2760 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#05#),
      2785 => to_slv(opcode_type, 16#01#),
      2786 => to_slv(opcode_type, 16#06#),
      2787 => to_slv(opcode_type, 16#09#),
      2788 => to_slv(opcode_type, 16#11#),
      2789 => to_slv(opcode_type, 16#0E#),
      2790 => to_slv(opcode_type, 16#02#),
      2791 => to_slv(opcode_type, 16#12#),
      2792 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#03#),
      2817 => to_slv(opcode_type, 16#05#),
      2818 => to_slv(opcode_type, 16#08#),
      2819 => to_slv(opcode_type, 16#04#),
      2820 => to_slv(opcode_type, 16#11#),
      2821 => to_slv(opcode_type, 16#07#),
      2822 => to_slv(opcode_type, 16#0C#),
      2823 => to_slv(opcode_type, 16#0D#),
      2824 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#04#),
      2849 => to_slv(opcode_type, 16#01#),
      2850 => to_slv(opcode_type, 16#06#),
      2851 => to_slv(opcode_type, 16#03#),
      2852 => to_slv(opcode_type, 16#0B#),
      2853 => to_slv(opcode_type, 16#08#),
      2854 => to_slv(opcode_type, 16#0A#),
      2855 => to_slv(opcode_type, 16#11#),
      2856 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#09#),
      2881 => to_slv(opcode_type, 16#09#),
      2882 => to_slv(opcode_type, 16#09#),
      2883 => to_slv(opcode_type, 16#01#),
      2884 => to_slv(opcode_type, 16#10#),
      2885 => to_slv(opcode_type, 16#0A#),
      2886 => to_slv(opcode_type, 16#0F#),
      2887 => to_slv(opcode_type, 16#11#),
      2888 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#02#),
      2913 => to_slv(opcode_type, 16#03#),
      2914 => to_slv(opcode_type, 16#09#),
      2915 => to_slv(opcode_type, 16#05#),
      2916 => to_slv(opcode_type, 16#0C#),
      2917 => to_slv(opcode_type, 16#06#),
      2918 => to_slv(opcode_type, 16#0F#),
      2919 => to_slv(opcode_type, 16#0B#),
      2920 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#05#),
      2945 => to_slv(opcode_type, 16#01#),
      2946 => to_slv(opcode_type, 16#09#),
      2947 => to_slv(opcode_type, 16#09#),
      2948 => to_slv(opcode_type, 16#0E#),
      2949 => to_slv(opcode_type, 16#0B#),
      2950 => to_slv(opcode_type, 16#03#),
      2951 => to_slv(opcode_type, 16#0F#),
      2952 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#09#),
      2977 => to_slv(opcode_type, 16#07#),
      2978 => to_slv(opcode_type, 16#05#),
      2979 => to_slv(opcode_type, 16#09#),
      2980 => to_slv(opcode_type, 16#0E#),
      2981 => to_slv(opcode_type, 16#0C#),
      2982 => to_slv(opcode_type, 16#0B#),
      2983 => to_slv(opcode_type, 16#0E#),
      2984 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#01#),
      3009 => to_slv(opcode_type, 16#05#),
      3010 => to_slv(opcode_type, 16#08#),
      3011 => to_slv(opcode_type, 16#04#),
      3012 => to_slv(opcode_type, 16#0D#),
      3013 => to_slv(opcode_type, 16#07#),
      3014 => to_slv(opcode_type, 16#0E#),
      3015 => to_slv(opcode_type, 16#A7#),
      3016 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#07#),
      3041 => to_slv(opcode_type, 16#07#),
      3042 => to_slv(opcode_type, 16#07#),
      3043 => to_slv(opcode_type, 16#05#),
      3044 => to_slv(opcode_type, 16#4C#),
      3045 => to_slv(opcode_type, 16#0C#),
      3046 => to_slv(opcode_type, 16#10#),
      3047 => to_slv(opcode_type, 16#38#),
      3048 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#07#),
      3073 => to_slv(opcode_type, 16#06#),
      3074 => to_slv(opcode_type, 16#08#),
      3075 => to_slv(opcode_type, 16#03#),
      3076 => to_slv(opcode_type, 16#0A#),
      3077 => to_slv(opcode_type, 16#0C#),
      3078 => to_slv(opcode_type, 16#0F#),
      3079 => to_slv(opcode_type, 16#11#),
      3080 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#03#),
      3105 => to_slv(opcode_type, 16#08#),
      3106 => to_slv(opcode_type, 16#08#),
      3107 => to_slv(opcode_type, 16#09#),
      3108 => to_slv(opcode_type, 16#0C#),
      3109 => to_slv(opcode_type, 16#0F#),
      3110 => to_slv(opcode_type, 16#0A#),
      3111 => to_slv(opcode_type, 16#10#),
      3112 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#05#),
      3137 => to_slv(opcode_type, 16#03#),
      3138 => to_slv(opcode_type, 16#08#),
      3139 => to_slv(opcode_type, 16#01#),
      3140 => to_slv(opcode_type, 16#0C#),
      3141 => to_slv(opcode_type, 16#06#),
      3142 => to_slv(opcode_type, 16#11#),
      3143 => to_slv(opcode_type, 16#0F#),
      3144 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#04#),
      3169 => to_slv(opcode_type, 16#08#),
      3170 => to_slv(opcode_type, 16#03#),
      3171 => to_slv(opcode_type, 16#01#),
      3172 => to_slv(opcode_type, 16#0E#),
      3173 => to_slv(opcode_type, 16#09#),
      3174 => to_slv(opcode_type, 16#0A#),
      3175 => to_slv(opcode_type, 16#0F#),
      3176 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#06#),
      3201 => to_slv(opcode_type, 16#07#),
      3202 => to_slv(opcode_type, 16#05#),
      3203 => to_slv(opcode_type, 16#03#),
      3204 => to_slv(opcode_type, 16#0C#),
      3205 => to_slv(opcode_type, 16#02#),
      3206 => to_slv(opcode_type, 16#10#),
      3207 => to_slv(opcode_type, 16#0C#),
      3208 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#01#),
      3234 => to_slv(opcode_type, 16#09#),
      3235 => to_slv(opcode_type, 16#07#),
      3236 => to_slv(opcode_type, 16#0C#),
      3237 => to_slv(opcode_type, 16#0A#),
      3238 => to_slv(opcode_type, 16#0A#),
      3239 => to_slv(opcode_type, 16#A9#),
      3240 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#03#),
      3265 => to_slv(opcode_type, 16#07#),
      3266 => to_slv(opcode_type, 16#08#),
      3267 => to_slv(opcode_type, 16#02#),
      3268 => to_slv(opcode_type, 16#0D#),
      3269 => to_slv(opcode_type, 16#03#),
      3270 => to_slv(opcode_type, 16#9D#),
      3271 => to_slv(opcode_type, 16#0D#),
      3272 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#09#),
      3297 => to_slv(opcode_type, 16#01#),
      3298 => to_slv(opcode_type, 16#05#),
      3299 => to_slv(opcode_type, 16#01#),
      3300 => to_slv(opcode_type, 16#0D#),
      3301 => to_slv(opcode_type, 16#08#),
      3302 => to_slv(opcode_type, 16#10#),
      3303 => to_slv(opcode_type, 16#10#),
      3304 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#01#),
      3329 => to_slv(opcode_type, 16#04#),
      3330 => to_slv(opcode_type, 16#09#),
      3331 => to_slv(opcode_type, 16#03#),
      3332 => to_slv(opcode_type, 16#0C#),
      3333 => to_slv(opcode_type, 16#06#),
      3334 => to_slv(opcode_type, 16#0C#),
      3335 => to_slv(opcode_type, 16#0B#),
      3336 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#09#),
      3361 => to_slv(opcode_type, 16#05#),
      3362 => to_slv(opcode_type, 16#01#),
      3363 => to_slv(opcode_type, 16#07#),
      3364 => to_slv(opcode_type, 16#0E#),
      3365 => to_slv(opcode_type, 16#0B#),
      3366 => to_slv(opcode_type, 16#04#),
      3367 => to_slv(opcode_type, 16#10#),
      3368 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#08#),
      3393 => to_slv(opcode_type, 16#06#),
      3394 => to_slv(opcode_type, 16#02#),
      3395 => to_slv(opcode_type, 16#01#),
      3396 => to_slv(opcode_type, 16#11#),
      3397 => to_slv(opcode_type, 16#04#),
      3398 => to_slv(opcode_type, 16#11#),
      3399 => to_slv(opcode_type, 16#0C#),
      3400 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#06#),
      3426 => to_slv(opcode_type, 16#01#),
      3427 => to_slv(opcode_type, 16#09#),
      3428 => to_slv(opcode_type, 16#0A#),
      3429 => to_slv(opcode_type, 16#0D#),
      3430 => to_slv(opcode_type, 16#11#),
      3431 => to_slv(opcode_type, 16#EE#),
      3432 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#03#),
      3457 => to_slv(opcode_type, 16#04#),
      3458 => to_slv(opcode_type, 16#08#),
      3459 => to_slv(opcode_type, 16#09#),
      3460 => to_slv(opcode_type, 16#B6#),
      3461 => to_slv(opcode_type, 16#11#),
      3462 => to_slv(opcode_type, 16#02#),
      3463 => to_slv(opcode_type, 16#0E#),
      3464 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#06#),
      3489 => to_slv(opcode_type, 16#06#),
      3490 => to_slv(opcode_type, 16#02#),
      3491 => to_slv(opcode_type, 16#08#),
      3492 => to_slv(opcode_type, 16#0B#),
      3493 => to_slv(opcode_type, 16#0B#),
      3494 => to_slv(opcode_type, 16#10#),
      3495 => to_slv(opcode_type, 16#0A#),
      3496 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#01#),
      3521 => to_slv(opcode_type, 16#07#),
      3522 => to_slv(opcode_type, 16#07#),
      3523 => to_slv(opcode_type, 16#07#),
      3524 => to_slv(opcode_type, 16#1C#),
      3525 => to_slv(opcode_type, 16#0C#),
      3526 => to_slv(opcode_type, 16#C5#),
      3527 => to_slv(opcode_type, 16#0C#),
      3528 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#08#),
      3553 => to_slv(opcode_type, 16#08#),
      3554 => to_slv(opcode_type, 16#01#),
      3555 => to_slv(opcode_type, 16#04#),
      3556 => to_slv(opcode_type, 16#0A#),
      3557 => to_slv(opcode_type, 16#04#),
      3558 => to_slv(opcode_type, 16#0C#),
      3559 => to_slv(opcode_type, 16#0E#),
      3560 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#02#),
      3585 => to_slv(opcode_type, 16#05#),
      3586 => to_slv(opcode_type, 16#07#),
      3587 => to_slv(opcode_type, 16#08#),
      3588 => to_slv(opcode_type, 16#0E#),
      3589 => to_slv(opcode_type, 16#10#),
      3590 => to_slv(opcode_type, 16#05#),
      3591 => to_slv(opcode_type, 16#0F#),
      3592 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#08#),
      3617 => to_slv(opcode_type, 16#03#),
      3618 => to_slv(opcode_type, 16#01#),
      3619 => to_slv(opcode_type, 16#01#),
      3620 => to_slv(opcode_type, 16#0B#),
      3621 => to_slv(opcode_type, 16#09#),
      3622 => to_slv(opcode_type, 16#11#),
      3623 => to_slv(opcode_type, 16#0A#),
      3624 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#06#),
      3649 => to_slv(opcode_type, 16#01#),
      3650 => to_slv(opcode_type, 16#03#),
      3651 => to_slv(opcode_type, 16#06#),
      3652 => to_slv(opcode_type, 16#0E#),
      3653 => to_slv(opcode_type, 16#0C#),
      3654 => to_slv(opcode_type, 16#05#),
      3655 => to_slv(opcode_type, 16#0B#),
      3656 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#02#),
      3681 => to_slv(opcode_type, 16#08#),
      3682 => to_slv(opcode_type, 16#06#),
      3683 => to_slv(opcode_type, 16#03#),
      3684 => to_slv(opcode_type, 16#0D#),
      3685 => to_slv(opcode_type, 16#01#),
      3686 => to_slv(opcode_type, 16#11#),
      3687 => to_slv(opcode_type, 16#0C#),
      3688 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#02#),
      3713 => to_slv(opcode_type, 16#01#),
      3714 => to_slv(opcode_type, 16#08#),
      3715 => to_slv(opcode_type, 16#06#),
      3716 => to_slv(opcode_type, 16#0D#),
      3717 => to_slv(opcode_type, 16#11#),
      3718 => to_slv(opcode_type, 16#01#),
      3719 => to_slv(opcode_type, 16#0B#),
      3720 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#03#),
      3745 => to_slv(opcode_type, 16#07#),
      3746 => to_slv(opcode_type, 16#06#),
      3747 => to_slv(opcode_type, 16#08#),
      3748 => to_slv(opcode_type, 16#0B#),
      3749 => to_slv(opcode_type, 16#0A#),
      3750 => to_slv(opcode_type, 16#0E#),
      3751 => to_slv(opcode_type, 16#0B#),
      3752 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#06#),
      3777 => to_slv(opcode_type, 16#04#),
      3778 => to_slv(opcode_type, 16#04#),
      3779 => to_slv(opcode_type, 16#06#),
      3780 => to_slv(opcode_type, 16#10#),
      3781 => to_slv(opcode_type, 16#10#),
      3782 => to_slv(opcode_type, 16#04#),
      3783 => to_slv(opcode_type, 16#E2#),
      3784 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#05#),
      3809 => to_slv(opcode_type, 16#03#),
      3810 => to_slv(opcode_type, 16#06#),
      3811 => to_slv(opcode_type, 16#01#),
      3812 => to_slv(opcode_type, 16#0F#),
      3813 => to_slv(opcode_type, 16#07#),
      3814 => to_slv(opcode_type, 16#11#),
      3815 => to_slv(opcode_type, 16#0A#),
      3816 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#04#),
      3841 => to_slv(opcode_type, 16#04#),
      3842 => to_slv(opcode_type, 16#06#),
      3843 => to_slv(opcode_type, 16#07#),
      3844 => to_slv(opcode_type, 16#10#),
      3845 => to_slv(opcode_type, 16#0D#),
      3846 => to_slv(opcode_type, 16#02#),
      3847 => to_slv(opcode_type, 16#0A#),
      3848 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#05#),
      3873 => to_slv(opcode_type, 16#05#),
      3874 => to_slv(opcode_type, 16#08#),
      3875 => to_slv(opcode_type, 16#06#),
      3876 => to_slv(opcode_type, 16#0C#),
      3877 => to_slv(opcode_type, 16#0C#),
      3878 => to_slv(opcode_type, 16#03#),
      3879 => to_slv(opcode_type, 16#11#),
      3880 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#02#),
      3905 => to_slv(opcode_type, 16#02#),
      3906 => to_slv(opcode_type, 16#07#),
      3907 => to_slv(opcode_type, 16#05#),
      3908 => to_slv(opcode_type, 16#10#),
      3909 => to_slv(opcode_type, 16#07#),
      3910 => to_slv(opcode_type, 16#11#),
      3911 => to_slv(opcode_type, 16#0F#),
      3912 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#09#),
      3937 => to_slv(opcode_type, 16#03#),
      3938 => to_slv(opcode_type, 16#06#),
      3939 => to_slv(opcode_type, 16#01#),
      3940 => to_slv(opcode_type, 16#0B#),
      3941 => to_slv(opcode_type, 16#03#),
      3942 => to_slv(opcode_type, 16#0B#),
      3943 => to_slv(opcode_type, 16#10#),
      3944 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#03#),
      3969 => to_slv(opcode_type, 16#08#),
      3970 => to_slv(opcode_type, 16#03#),
      3971 => to_slv(opcode_type, 16#05#),
      3972 => to_slv(opcode_type, 16#0F#),
      3973 => to_slv(opcode_type, 16#05#),
      3974 => to_slv(opcode_type, 16#03#),
      3975 => to_slv(opcode_type, 16#11#),
      3976 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#09#),
      4001 => to_slv(opcode_type, 16#09#),
      4002 => to_slv(opcode_type, 16#07#),
      4003 => to_slv(opcode_type, 16#01#),
      4004 => to_slv(opcode_type, 16#10#),
      4005 => to_slv(opcode_type, 16#0B#),
      4006 => to_slv(opcode_type, 16#0C#),
      4007 => to_slv(opcode_type, 16#10#),
      4008 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#02#),
      4033 => to_slv(opcode_type, 16#09#),
      4034 => to_slv(opcode_type, 16#01#),
      4035 => to_slv(opcode_type, 16#02#),
      4036 => to_slv(opcode_type, 16#0B#),
      4037 => to_slv(opcode_type, 16#05#),
      4038 => to_slv(opcode_type, 16#04#),
      4039 => to_slv(opcode_type, 16#0D#),
      4040 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#08#),
      4065 => to_slv(opcode_type, 16#01#),
      4066 => to_slv(opcode_type, 16#04#),
      4067 => to_slv(opcode_type, 16#03#),
      4068 => to_slv(opcode_type, 16#0A#),
      4069 => to_slv(opcode_type, 16#09#),
      4070 => to_slv(opcode_type, 16#0E#),
      4071 => to_slv(opcode_type, 16#11#),
      4072 to 4095 => (others => '0')
  ),

    -- Bin `9`...
    8 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#04#),
      1 => to_slv(opcode_type, 16#02#),
      2 => to_slv(opcode_type, 16#06#),
      3 => to_slv(opcode_type, 16#08#),
      4 => to_slv(opcode_type, 16#0A#),
      5 => to_slv(opcode_type, 16#10#),
      6 => to_slv(opcode_type, 16#09#),
      7 => to_slv(opcode_type, 16#FD#),
      8 => to_slv(opcode_type, 16#0C#),
      9 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#03#),
      33 => to_slv(opcode_type, 16#03#),
      34 => to_slv(opcode_type, 16#09#),
      35 => to_slv(opcode_type, 16#07#),
      36 => to_slv(opcode_type, 16#10#),
      37 => to_slv(opcode_type, 16#78#),
      38 => to_slv(opcode_type, 16#06#),
      39 => to_slv(opcode_type, 16#0E#),
      40 => to_slv(opcode_type, 16#11#),
      41 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#03#),
      65 => to_slv(opcode_type, 16#02#),
      66 => to_slv(opcode_type, 16#07#),
      67 => to_slv(opcode_type, 16#06#),
      68 => to_slv(opcode_type, 16#0E#),
      69 => to_slv(opcode_type, 16#10#),
      70 => to_slv(opcode_type, 16#06#),
      71 => to_slv(opcode_type, 16#11#),
      72 => to_slv(opcode_type, 16#0E#),
      73 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#08#),
      97 => to_slv(opcode_type, 16#04#),
      98 => to_slv(opcode_type, 16#05#),
      99 => to_slv(opcode_type, 16#03#),
      100 => to_slv(opcode_type, 16#0A#),
      101 => to_slv(opcode_type, 16#02#),
      102 => to_slv(opcode_type, 16#08#),
      103 => to_slv(opcode_type, 16#11#),
      104 => to_slv(opcode_type, 16#0D#),
      105 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#03#),
      129 => to_slv(opcode_type, 16#09#),
      130 => to_slv(opcode_type, 16#07#),
      131 => to_slv(opcode_type, 16#07#),
      132 => to_slv(opcode_type, 16#11#),
      133 => to_slv(opcode_type, 16#0E#),
      134 => to_slv(opcode_type, 16#05#),
      135 => to_slv(opcode_type, 16#11#),
      136 => to_slv(opcode_type, 16#80#),
      137 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#06#),
      161 => to_slv(opcode_type, 16#09#),
      162 => to_slv(opcode_type, 16#02#),
      163 => to_slv(opcode_type, 16#09#),
      164 => to_slv(opcode_type, 16#80#),
      165 => to_slv(opcode_type, 16#10#),
      166 => to_slv(opcode_type, 16#04#),
      167 => to_slv(opcode_type, 16#0C#),
      168 => to_slv(opcode_type, 16#11#),
      169 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#03#),
      193 => to_slv(opcode_type, 16#09#),
      194 => to_slv(opcode_type, 16#01#),
      195 => to_slv(opcode_type, 16#04#),
      196 => to_slv(opcode_type, 16#10#),
      197 => to_slv(opcode_type, 16#06#),
      198 => to_slv(opcode_type, 16#02#),
      199 => to_slv(opcode_type, 16#0B#),
      200 => to_slv(opcode_type, 16#0D#),
      201 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#01#),
      225 => to_slv(opcode_type, 16#01#),
      226 => to_slv(opcode_type, 16#07#),
      227 => to_slv(opcode_type, 16#06#),
      228 => to_slv(opcode_type, 16#0A#),
      229 => to_slv(opcode_type, 16#0A#),
      230 => to_slv(opcode_type, 16#09#),
      231 => to_slv(opcode_type, 16#0B#),
      232 => to_slv(opcode_type, 16#0A#),
      233 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#07#),
      257 => to_slv(opcode_type, 16#08#),
      258 => to_slv(opcode_type, 16#03#),
      259 => to_slv(opcode_type, 16#03#),
      260 => to_slv(opcode_type, 16#0D#),
      261 => to_slv(opcode_type, 16#05#),
      262 => to_slv(opcode_type, 16#01#),
      263 => to_slv(opcode_type, 16#0A#),
      264 => to_slv(opcode_type, 16#0E#),
      265 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#05#),
      289 => to_slv(opcode_type, 16#07#),
      290 => to_slv(opcode_type, 16#02#),
      291 => to_slv(opcode_type, 16#02#),
      292 => to_slv(opcode_type, 16#0C#),
      293 => to_slv(opcode_type, 16#09#),
      294 => to_slv(opcode_type, 16#02#),
      295 => to_slv(opcode_type, 16#6C#),
      296 => to_slv(opcode_type, 16#0E#),
      297 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#08#),
      321 => to_slv(opcode_type, 16#03#),
      322 => to_slv(opcode_type, 16#06#),
      323 => to_slv(opcode_type, 16#03#),
      324 => to_slv(opcode_type, 16#0A#),
      325 => to_slv(opcode_type, 16#01#),
      326 => to_slv(opcode_type, 16#BF#),
      327 => to_slv(opcode_type, 16#02#),
      328 => to_slv(opcode_type, 16#0A#),
      329 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#03#),
      353 => to_slv(opcode_type, 16#03#),
      354 => to_slv(opcode_type, 16#07#),
      355 => to_slv(opcode_type, 16#08#),
      356 => to_slv(opcode_type, 16#10#),
      357 => to_slv(opcode_type, 16#67#),
      358 => to_slv(opcode_type, 16#07#),
      359 => to_slv(opcode_type, 16#0A#),
      360 => to_slv(opcode_type, 16#10#),
      361 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#09#),
      385 => to_slv(opcode_type, 16#03#),
      386 => to_slv(opcode_type, 16#09#),
      387 => to_slv(opcode_type, 16#06#),
      388 => to_slv(opcode_type, 16#0E#),
      389 => to_slv(opcode_type, 16#10#),
      390 => to_slv(opcode_type, 16#01#),
      391 => to_slv(opcode_type, 16#0F#),
      392 => to_slv(opcode_type, 16#0A#),
      393 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#07#),
      417 => to_slv(opcode_type, 16#01#),
      418 => to_slv(opcode_type, 16#08#),
      419 => to_slv(opcode_type, 16#02#),
      420 => to_slv(opcode_type, 16#0F#),
      421 => to_slv(opcode_type, 16#07#),
      422 => to_slv(opcode_type, 16#10#),
      423 => to_slv(opcode_type, 16#0F#),
      424 => to_slv(opcode_type, 16#10#),
      425 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#04#),
      449 => to_slv(opcode_type, 16#07#),
      450 => to_slv(opcode_type, 16#01#),
      451 => to_slv(opcode_type, 16#06#),
      452 => to_slv(opcode_type, 16#11#),
      453 => to_slv(opcode_type, 16#0C#),
      454 => to_slv(opcode_type, 16#03#),
      455 => to_slv(opcode_type, 16#04#),
      456 => to_slv(opcode_type, 16#0A#),
      457 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#04#),
      481 => to_slv(opcode_type, 16#03#),
      482 => to_slv(opcode_type, 16#08#),
      483 => to_slv(opcode_type, 16#08#),
      484 => to_slv(opcode_type, 16#0B#),
      485 => to_slv(opcode_type, 16#0C#),
      486 => to_slv(opcode_type, 16#07#),
      487 => to_slv(opcode_type, 16#11#),
      488 => to_slv(opcode_type, 16#0E#),
      489 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#01#),
      513 => to_slv(opcode_type, 16#03#),
      514 => to_slv(opcode_type, 16#07#),
      515 => to_slv(opcode_type, 16#08#),
      516 => to_slv(opcode_type, 16#0D#),
      517 => to_slv(opcode_type, 16#0A#),
      518 => to_slv(opcode_type, 16#07#),
      519 => to_slv(opcode_type, 16#0A#),
      520 => to_slv(opcode_type, 16#10#),
      521 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#05#),
      545 => to_slv(opcode_type, 16#01#),
      546 => to_slv(opcode_type, 16#07#),
      547 => to_slv(opcode_type, 16#08#),
      548 => to_slv(opcode_type, 16#0B#),
      549 => to_slv(opcode_type, 16#0B#),
      550 => to_slv(opcode_type, 16#07#),
      551 => to_slv(opcode_type, 16#0C#),
      552 => to_slv(opcode_type, 16#0E#),
      553 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#06#),
      577 => to_slv(opcode_type, 16#06#),
      578 => to_slv(opcode_type, 16#08#),
      579 => to_slv(opcode_type, 16#06#),
      580 => to_slv(opcode_type, 16#68#),
      581 => to_slv(opcode_type, 16#11#),
      582 => to_slv(opcode_type, 16#0B#),
      583 => to_slv(opcode_type, 16#0F#),
      584 => to_slv(opcode_type, 16#10#),
      585 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#04#),
      609 => to_slv(opcode_type, 16#08#),
      610 => to_slv(opcode_type, 16#09#),
      611 => to_slv(opcode_type, 16#01#),
      612 => to_slv(opcode_type, 16#0C#),
      613 => to_slv(opcode_type, 16#08#),
      614 => to_slv(opcode_type, 16#0D#),
      615 => to_slv(opcode_type, 16#0A#),
      616 => to_slv(opcode_type, 16#0C#),
      617 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#02#),
      641 => to_slv(opcode_type, 16#03#),
      642 => to_slv(opcode_type, 16#08#),
      643 => to_slv(opcode_type, 16#07#),
      644 => to_slv(opcode_type, 16#0D#),
      645 => to_slv(opcode_type, 16#10#),
      646 => to_slv(opcode_type, 16#09#),
      647 => to_slv(opcode_type, 16#4F#),
      648 => to_slv(opcode_type, 16#0A#),
      649 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#08#),
      673 => to_slv(opcode_type, 16#04#),
      674 => to_slv(opcode_type, 16#08#),
      675 => to_slv(opcode_type, 16#08#),
      676 => to_slv(opcode_type, 16#0E#),
      677 => to_slv(opcode_type, 16#CB#),
      678 => to_slv(opcode_type, 16#01#),
      679 => to_slv(opcode_type, 16#0D#),
      680 => to_slv(opcode_type, 16#8E#),
      681 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#04#),
      705 => to_slv(opcode_type, 16#09#),
      706 => to_slv(opcode_type, 16#05#),
      707 => to_slv(opcode_type, 16#06#),
      708 => to_slv(opcode_type, 16#11#),
      709 => to_slv(opcode_type, 16#30#),
      710 => to_slv(opcode_type, 16#08#),
      711 => to_slv(opcode_type, 16#0C#),
      712 => to_slv(opcode_type, 16#0E#),
      713 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#04#),
      737 => to_slv(opcode_type, 16#06#),
      738 => to_slv(opcode_type, 16#01#),
      739 => to_slv(opcode_type, 16#06#),
      740 => to_slv(opcode_type, 16#11#),
      741 => to_slv(opcode_type, 16#62#),
      742 => to_slv(opcode_type, 16#07#),
      743 => to_slv(opcode_type, 16#0E#),
      744 => to_slv(opcode_type, 16#11#),
      745 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#05#),
      769 => to_slv(opcode_type, 16#06#),
      770 => to_slv(opcode_type, 16#05#),
      771 => to_slv(opcode_type, 16#05#),
      772 => to_slv(opcode_type, 16#0F#),
      773 => to_slv(opcode_type, 16#05#),
      774 => to_slv(opcode_type, 16#08#),
      775 => to_slv(opcode_type, 16#0D#),
      776 => to_slv(opcode_type, 16#0E#),
      777 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#02#),
      801 => to_slv(opcode_type, 16#07#),
      802 => to_slv(opcode_type, 16#01#),
      803 => to_slv(opcode_type, 16#03#),
      804 => to_slv(opcode_type, 16#10#),
      805 => to_slv(opcode_type, 16#03#),
      806 => to_slv(opcode_type, 16#07#),
      807 => to_slv(opcode_type, 16#10#),
      808 => to_slv(opcode_type, 16#0D#),
      809 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#06#),
      833 => to_slv(opcode_type, 16#04#),
      834 => to_slv(opcode_type, 16#01#),
      835 => to_slv(opcode_type, 16#08#),
      836 => to_slv(opcode_type, 16#0F#),
      837 => to_slv(opcode_type, 16#11#),
      838 => to_slv(opcode_type, 16#08#),
      839 => to_slv(opcode_type, 16#0F#),
      840 => to_slv(opcode_type, 16#0C#),
      841 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#09#),
      865 => to_slv(opcode_type, 16#01#),
      866 => to_slv(opcode_type, 16#03#),
      867 => to_slv(opcode_type, 16#02#),
      868 => to_slv(opcode_type, 16#10#),
      869 => to_slv(opcode_type, 16#06#),
      870 => to_slv(opcode_type, 16#01#),
      871 => to_slv(opcode_type, 16#0C#),
      872 => to_slv(opcode_type, 16#0B#),
      873 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#06#),
      898 => to_slv(opcode_type, 16#04#),
      899 => to_slv(opcode_type, 16#04#),
      900 => to_slv(opcode_type, 16#0E#),
      901 => to_slv(opcode_type, 16#06#),
      902 => to_slv(opcode_type, 16#0C#),
      903 => to_slv(opcode_type, 16#0C#),
      904 => to_slv(opcode_type, 16#3E#),
      905 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#03#),
      929 => to_slv(opcode_type, 16#08#),
      930 => to_slv(opcode_type, 16#07#),
      931 => to_slv(opcode_type, 16#06#),
      932 => to_slv(opcode_type, 16#32#),
      933 => to_slv(opcode_type, 16#D4#),
      934 => to_slv(opcode_type, 16#03#),
      935 => to_slv(opcode_type, 16#0D#),
      936 => to_slv(opcode_type, 16#10#),
      937 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#01#),
      961 => to_slv(opcode_type, 16#05#),
      962 => to_slv(opcode_type, 16#09#),
      963 => to_slv(opcode_type, 16#06#),
      964 => to_slv(opcode_type, 16#11#),
      965 => to_slv(opcode_type, 16#0D#),
      966 => to_slv(opcode_type, 16#06#),
      967 => to_slv(opcode_type, 16#0A#),
      968 => to_slv(opcode_type, 16#11#),
      969 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#04#),
      993 => to_slv(opcode_type, 16#04#),
      994 => to_slv(opcode_type, 16#08#),
      995 => to_slv(opcode_type, 16#06#),
      996 => to_slv(opcode_type, 16#0F#),
      997 => to_slv(opcode_type, 16#0B#),
      998 => to_slv(opcode_type, 16#08#),
      999 => to_slv(opcode_type, 16#0A#),
      1000 => to_slv(opcode_type, 16#0F#),
      1001 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#09#),
      1025 => to_slv(opcode_type, 16#07#),
      1026 => to_slv(opcode_type, 16#06#),
      1027 => to_slv(opcode_type, 16#06#),
      1028 => to_slv(opcode_type, 16#67#),
      1029 => to_slv(opcode_type, 16#10#),
      1030 => to_slv(opcode_type, 16#0D#),
      1031 => to_slv(opcode_type, 16#10#),
      1032 => to_slv(opcode_type, 16#11#),
      1033 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#04#),
      1057 => to_slv(opcode_type, 16#06#),
      1058 => to_slv(opcode_type, 16#01#),
      1059 => to_slv(opcode_type, 16#06#),
      1060 => to_slv(opcode_type, 16#0D#),
      1061 => to_slv(opcode_type, 16#6A#),
      1062 => to_slv(opcode_type, 16#06#),
      1063 => to_slv(opcode_type, 16#0B#),
      1064 => to_slv(opcode_type, 16#0F#),
      1065 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#03#),
      1089 => to_slv(opcode_type, 16#09#),
      1090 => to_slv(opcode_type, 16#09#),
      1091 => to_slv(opcode_type, 16#01#),
      1092 => to_slv(opcode_type, 16#0E#),
      1093 => to_slv(opcode_type, 16#09#),
      1094 => to_slv(opcode_type, 16#0A#),
      1095 => to_slv(opcode_type, 16#10#),
      1096 => to_slv(opcode_type, 16#0D#),
      1097 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#03#),
      1121 => to_slv(opcode_type, 16#04#),
      1122 => to_slv(opcode_type, 16#09#),
      1123 => to_slv(opcode_type, 16#09#),
      1124 => to_slv(opcode_type, 16#0C#),
      1125 => to_slv(opcode_type, 16#8D#),
      1126 => to_slv(opcode_type, 16#07#),
      1127 => to_slv(opcode_type, 16#0C#),
      1128 => to_slv(opcode_type, 16#FD#),
      1129 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#06#),
      1153 => to_slv(opcode_type, 16#07#),
      1154 => to_slv(opcode_type, 16#02#),
      1155 => to_slv(opcode_type, 16#07#),
      1156 => to_slv(opcode_type, 16#0F#),
      1157 => to_slv(opcode_type, 16#0B#),
      1158 => to_slv(opcode_type, 16#02#),
      1159 => to_slv(opcode_type, 16#10#),
      1160 => to_slv(opcode_type, 16#0E#),
      1161 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#07#),
      1185 => to_slv(opcode_type, 16#08#),
      1186 => to_slv(opcode_type, 16#01#),
      1187 => to_slv(opcode_type, 16#04#),
      1188 => to_slv(opcode_type, 16#11#),
      1189 => to_slv(opcode_type, 16#07#),
      1190 => to_slv(opcode_type, 16#11#),
      1191 => to_slv(opcode_type, 16#11#),
      1192 => to_slv(opcode_type, 16#45#),
      1193 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#07#),
      1217 => to_slv(opcode_type, 16#06#),
      1218 => to_slv(opcode_type, 16#02#),
      1219 => to_slv(opcode_type, 16#05#),
      1220 => to_slv(opcode_type, 16#10#),
      1221 => to_slv(opcode_type, 16#09#),
      1222 => to_slv(opcode_type, 16#5E#),
      1223 => to_slv(opcode_type, 16#11#),
      1224 => to_slv(opcode_type, 16#0F#),
      1225 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#05#),
      1249 => to_slv(opcode_type, 16#09#),
      1250 => to_slv(opcode_type, 16#07#),
      1251 => to_slv(opcode_type, 16#07#),
      1252 => to_slv(opcode_type, 16#0E#),
      1253 => to_slv(opcode_type, 16#0A#),
      1254 => to_slv(opcode_type, 16#04#),
      1255 => to_slv(opcode_type, 16#0F#),
      1256 => to_slv(opcode_type, 16#79#),
      1257 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#07#),
      1282 => to_slv(opcode_type, 16#07#),
      1283 => to_slv(opcode_type, 16#04#),
      1284 => to_slv(opcode_type, 16#0B#),
      1285 => to_slv(opcode_type, 16#01#),
      1286 => to_slv(opcode_type, 16#11#),
      1287 => to_slv(opcode_type, 16#0C#),
      1288 => to_slv(opcode_type, 16#0E#),
      1289 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#07#),
      1313 => to_slv(opcode_type, 16#05#),
      1314 => to_slv(opcode_type, 16#05#),
      1315 => to_slv(opcode_type, 16#09#),
      1316 => to_slv(opcode_type, 16#0F#),
      1317 => to_slv(opcode_type, 16#B0#),
      1318 => to_slv(opcode_type, 16#08#),
      1319 => to_slv(opcode_type, 16#0B#),
      1320 => to_slv(opcode_type, 16#0B#),
      1321 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#03#),
      1345 => to_slv(opcode_type, 16#09#),
      1346 => to_slv(opcode_type, 16#06#),
      1347 => to_slv(opcode_type, 16#07#),
      1348 => to_slv(opcode_type, 16#6F#),
      1349 => to_slv(opcode_type, 16#11#),
      1350 => to_slv(opcode_type, 16#04#),
      1351 => to_slv(opcode_type, 16#10#),
      1352 => to_slv(opcode_type, 16#11#),
      1353 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#02#),
      1377 => to_slv(opcode_type, 16#04#),
      1378 => to_slv(opcode_type, 16#07#),
      1379 => to_slv(opcode_type, 16#06#),
      1380 => to_slv(opcode_type, 16#0B#),
      1381 => to_slv(opcode_type, 16#0F#),
      1382 => to_slv(opcode_type, 16#06#),
      1383 => to_slv(opcode_type, 16#1D#),
      1384 => to_slv(opcode_type, 16#0E#),
      1385 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#08#),
      1409 => to_slv(opcode_type, 16#09#),
      1410 => to_slv(opcode_type, 16#02#),
      1411 => to_slv(opcode_type, 16#02#),
      1412 => to_slv(opcode_type, 16#0A#),
      1413 => to_slv(opcode_type, 16#09#),
      1414 => to_slv(opcode_type, 16#0D#),
      1415 => to_slv(opcode_type, 16#10#),
      1416 => to_slv(opcode_type, 16#0B#),
      1417 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#05#),
      1441 => to_slv(opcode_type, 16#06#),
      1442 => to_slv(opcode_type, 16#07#),
      1443 => to_slv(opcode_type, 16#08#),
      1444 => to_slv(opcode_type, 16#0F#),
      1445 => to_slv(opcode_type, 16#0B#),
      1446 => to_slv(opcode_type, 16#01#),
      1447 => to_slv(opcode_type, 16#0B#),
      1448 => to_slv(opcode_type, 16#0E#),
      1449 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#08#),
      1473 => to_slv(opcode_type, 16#09#),
      1474 => to_slv(opcode_type, 16#06#),
      1475 => to_slv(opcode_type, 16#06#),
      1476 => to_slv(opcode_type, 16#0C#),
      1477 => to_slv(opcode_type, 16#0B#),
      1478 => to_slv(opcode_type, 16#0F#),
      1479 => to_slv(opcode_type, 16#0F#),
      1480 => to_slv(opcode_type, 16#0F#),
      1481 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#07#),
      1505 => to_slv(opcode_type, 16#05#),
      1506 => to_slv(opcode_type, 16#03#),
      1507 => to_slv(opcode_type, 16#08#),
      1508 => to_slv(opcode_type, 16#0C#),
      1509 => to_slv(opcode_type, 16#11#),
      1510 => to_slv(opcode_type, 16#01#),
      1511 => to_slv(opcode_type, 16#03#),
      1512 => to_slv(opcode_type, 16#0F#),
      1513 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#07#),
      1537 => to_slv(opcode_type, 16#01#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#02#),
      1540 => to_slv(opcode_type, 16#0F#),
      1541 => to_slv(opcode_type, 16#09#),
      1542 => to_slv(opcode_type, 16#11#),
      1543 => to_slv(opcode_type, 16#11#),
      1544 => to_slv(opcode_type, 16#E9#),
      1545 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#06#),
      1569 => to_slv(opcode_type, 16#02#),
      1570 => to_slv(opcode_type, 16#07#),
      1571 => to_slv(opcode_type, 16#05#),
      1572 => to_slv(opcode_type, 16#0A#),
      1573 => to_slv(opcode_type, 16#03#),
      1574 => to_slv(opcode_type, 16#0E#),
      1575 => to_slv(opcode_type, 16#04#),
      1576 => to_slv(opcode_type, 16#0F#),
      1577 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#08#),
      1602 => to_slv(opcode_type, 16#02#),
      1603 => to_slv(opcode_type, 16#06#),
      1604 => to_slv(opcode_type, 16#97#),
      1605 => to_slv(opcode_type, 16#95#),
      1606 => to_slv(opcode_type, 16#04#),
      1607 => to_slv(opcode_type, 16#30#),
      1608 => to_slv(opcode_type, 16#95#),
      1609 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#04#),
      1633 => to_slv(opcode_type, 16#05#),
      1634 => to_slv(opcode_type, 16#07#),
      1635 => to_slv(opcode_type, 16#07#),
      1636 => to_slv(opcode_type, 16#0E#),
      1637 => to_slv(opcode_type, 16#0B#),
      1638 => to_slv(opcode_type, 16#08#),
      1639 => to_slv(opcode_type, 16#0C#),
      1640 => to_slv(opcode_type, 16#11#),
      1641 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#02#),
      1665 => to_slv(opcode_type, 16#04#),
      1666 => to_slv(opcode_type, 16#08#),
      1667 => to_slv(opcode_type, 16#08#),
      1668 => to_slv(opcode_type, 16#10#),
      1669 => to_slv(opcode_type, 16#10#),
      1670 => to_slv(opcode_type, 16#08#),
      1671 => to_slv(opcode_type, 16#50#),
      1672 => to_slv(opcode_type, 16#0D#),
      1673 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#08#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#08#),
      1699 => to_slv(opcode_type, 16#09#),
      1700 => to_slv(opcode_type, 16#95#),
      1701 => to_slv(opcode_type, 16#0C#),
      1702 => to_slv(opcode_type, 16#0D#),
      1703 => to_slv(opcode_type, 16#0E#),
      1704 => to_slv(opcode_type, 16#0C#),
      1705 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#09#),
      1729 => to_slv(opcode_type, 16#04#),
      1730 => to_slv(opcode_type, 16#03#),
      1731 => to_slv(opcode_type, 16#06#),
      1732 => to_slv(opcode_type, 16#0C#),
      1733 => to_slv(opcode_type, 16#0B#),
      1734 => to_slv(opcode_type, 16#01#),
      1735 => to_slv(opcode_type, 16#03#),
      1736 => to_slv(opcode_type, 16#0B#),
      1737 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#06#),
      1761 => to_slv(opcode_type, 16#01#),
      1762 => to_slv(opcode_type, 16#02#),
      1763 => to_slv(opcode_type, 16#03#),
      1764 => to_slv(opcode_type, 16#0D#),
      1765 => to_slv(opcode_type, 16#03#),
      1766 => to_slv(opcode_type, 16#04#),
      1767 => to_slv(opcode_type, 16#04#),
      1768 => to_slv(opcode_type, 16#0F#),
      1769 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#02#),
      1793 => to_slv(opcode_type, 16#01#),
      1794 => to_slv(opcode_type, 16#08#),
      1795 => to_slv(opcode_type, 16#09#),
      1796 => to_slv(opcode_type, 16#0C#),
      1797 => to_slv(opcode_type, 16#0D#),
      1798 => to_slv(opcode_type, 16#09#),
      1799 => to_slv(opcode_type, 16#0A#),
      1800 => to_slv(opcode_type, 16#0A#),
      1801 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#01#),
      1825 => to_slv(opcode_type, 16#04#),
      1826 => to_slv(opcode_type, 16#08#),
      1827 => to_slv(opcode_type, 16#06#),
      1828 => to_slv(opcode_type, 16#0D#),
      1829 => to_slv(opcode_type, 16#0C#),
      1830 => to_slv(opcode_type, 16#06#),
      1831 => to_slv(opcode_type, 16#0F#),
      1832 => to_slv(opcode_type, 16#0D#),
      1833 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#07#),
      1857 => to_slv(opcode_type, 16#09#),
      1858 => to_slv(opcode_type, 16#01#),
      1859 => to_slv(opcode_type, 16#04#),
      1860 => to_slv(opcode_type, 16#10#),
      1861 => to_slv(opcode_type, 16#08#),
      1862 => to_slv(opcode_type, 16#0D#),
      1863 => to_slv(opcode_type, 16#0D#),
      1864 => to_slv(opcode_type, 16#0F#),
      1865 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#05#),
      1889 => to_slv(opcode_type, 16#04#),
      1890 => to_slv(opcode_type, 16#06#),
      1891 => to_slv(opcode_type, 16#08#),
      1892 => to_slv(opcode_type, 16#0E#),
      1893 => to_slv(opcode_type, 16#0B#),
      1894 => to_slv(opcode_type, 16#08#),
      1895 => to_slv(opcode_type, 16#0C#),
      1896 => to_slv(opcode_type, 16#0A#),
      1897 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#02#),
      1921 => to_slv(opcode_type, 16#04#),
      1922 => to_slv(opcode_type, 16#08#),
      1923 => to_slv(opcode_type, 16#07#),
      1924 => to_slv(opcode_type, 16#0E#),
      1925 => to_slv(opcode_type, 16#0E#),
      1926 => to_slv(opcode_type, 16#09#),
      1927 => to_slv(opcode_type, 16#11#),
      1928 => to_slv(opcode_type, 16#11#),
      1929 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#01#),
      1953 => to_slv(opcode_type, 16#07#),
      1954 => to_slv(opcode_type, 16#01#),
      1955 => to_slv(opcode_type, 16#06#),
      1956 => to_slv(opcode_type, 16#0F#),
      1957 => to_slv(opcode_type, 16#11#),
      1958 => to_slv(opcode_type, 16#07#),
      1959 => to_slv(opcode_type, 16#0E#),
      1960 => to_slv(opcode_type, 16#10#),
      1961 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#05#),
      1985 => to_slv(opcode_type, 16#05#),
      1986 => to_slv(opcode_type, 16#08#),
      1987 => to_slv(opcode_type, 16#06#),
      1988 => to_slv(opcode_type, 16#0B#),
      1989 => to_slv(opcode_type, 16#10#),
      1990 => to_slv(opcode_type, 16#06#),
      1991 => to_slv(opcode_type, 16#0B#),
      1992 => to_slv(opcode_type, 16#20#),
      1993 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#03#),
      2017 => to_slv(opcode_type, 16#01#),
      2018 => to_slv(opcode_type, 16#06#),
      2019 => to_slv(opcode_type, 16#07#),
      2020 => to_slv(opcode_type, 16#11#),
      2021 => to_slv(opcode_type, 16#0A#),
      2022 => to_slv(opcode_type, 16#06#),
      2023 => to_slv(opcode_type, 16#10#),
      2024 => to_slv(opcode_type, 16#0E#),
      2025 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#06#),
      2049 => to_slv(opcode_type, 16#08#),
      2050 => to_slv(opcode_type, 16#09#),
      2051 => to_slv(opcode_type, 16#06#),
      2052 => to_slv(opcode_type, 16#0D#),
      2053 => to_slv(opcode_type, 16#9C#),
      2054 => to_slv(opcode_type, 16#11#),
      2055 => to_slv(opcode_type, 16#0E#),
      2056 => to_slv(opcode_type, 16#11#),
      2057 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#04#),
      2081 => to_slv(opcode_type, 16#08#),
      2082 => to_slv(opcode_type, 16#07#),
      2083 => to_slv(opcode_type, 16#02#),
      2084 => to_slv(opcode_type, 16#0C#),
      2085 => to_slv(opcode_type, 16#06#),
      2086 => to_slv(opcode_type, 16#0C#),
      2087 => to_slv(opcode_type, 16#2C#),
      2088 => to_slv(opcode_type, 16#11#),
      2089 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#01#),
      2113 => to_slv(opcode_type, 16#09#),
      2114 => to_slv(opcode_type, 16#01#),
      2115 => to_slv(opcode_type, 16#06#),
      2116 => to_slv(opcode_type, 16#0C#),
      2117 => to_slv(opcode_type, 16#0E#),
      2118 => to_slv(opcode_type, 16#02#),
      2119 => to_slv(opcode_type, 16#01#),
      2120 => to_slv(opcode_type, 16#0F#),
      2121 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#04#),
      2145 => to_slv(opcode_type, 16#04#),
      2146 => to_slv(opcode_type, 16#08#),
      2147 => to_slv(opcode_type, 16#06#),
      2148 => to_slv(opcode_type, 16#0C#),
      2149 => to_slv(opcode_type, 16#23#),
      2150 => to_slv(opcode_type, 16#07#),
      2151 => to_slv(opcode_type, 16#11#),
      2152 => to_slv(opcode_type, 16#0D#),
      2153 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#03#),
      2177 => to_slv(opcode_type, 16#01#),
      2178 => to_slv(opcode_type, 16#06#),
      2179 => to_slv(opcode_type, 16#06#),
      2180 => to_slv(opcode_type, 16#0C#),
      2181 => to_slv(opcode_type, 16#10#),
      2182 => to_slv(opcode_type, 16#09#),
      2183 => to_slv(opcode_type, 16#11#),
      2184 => to_slv(opcode_type, 16#0C#),
      2185 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#05#),
      2209 => to_slv(opcode_type, 16#04#),
      2210 => to_slv(opcode_type, 16#07#),
      2211 => to_slv(opcode_type, 16#07#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#10#),
      2214 => to_slv(opcode_type, 16#07#),
      2215 => to_slv(opcode_type, 16#0A#),
      2216 => to_slv(opcode_type, 16#10#),
      2217 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#04#),
      2241 => to_slv(opcode_type, 16#04#),
      2242 => to_slv(opcode_type, 16#08#),
      2243 => to_slv(opcode_type, 16#06#),
      2244 => to_slv(opcode_type, 16#0D#),
      2245 => to_slv(opcode_type, 16#0D#),
      2246 => to_slv(opcode_type, 16#08#),
      2247 => to_slv(opcode_type, 16#0D#),
      2248 => to_slv(opcode_type, 16#0F#),
      2249 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#02#),
      2273 => to_slv(opcode_type, 16#04#),
      2274 => to_slv(opcode_type, 16#06#),
      2275 => to_slv(opcode_type, 16#07#),
      2276 => to_slv(opcode_type, 16#0A#),
      2277 => to_slv(opcode_type, 16#0F#),
      2278 => to_slv(opcode_type, 16#06#),
      2279 => to_slv(opcode_type, 16#0D#),
      2280 => to_slv(opcode_type, 16#11#),
      2281 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#02#),
      2305 => to_slv(opcode_type, 16#08#),
      2306 => to_slv(opcode_type, 16#06#),
      2307 => to_slv(opcode_type, 16#01#),
      2308 => to_slv(opcode_type, 16#0A#),
      2309 => to_slv(opcode_type, 16#08#),
      2310 => to_slv(opcode_type, 16#0F#),
      2311 => to_slv(opcode_type, 16#E5#),
      2312 => to_slv(opcode_type, 16#0A#),
      2313 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#09#),
      2337 => to_slv(opcode_type, 16#08#),
      2338 => to_slv(opcode_type, 16#04#),
      2339 => to_slv(opcode_type, 16#01#),
      2340 => to_slv(opcode_type, 16#0C#),
      2341 => to_slv(opcode_type, 16#03#),
      2342 => to_slv(opcode_type, 16#01#),
      2343 => to_slv(opcode_type, 16#F8#),
      2344 => to_slv(opcode_type, 16#11#),
      2345 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#06#),
      2369 => to_slv(opcode_type, 16#01#),
      2370 => to_slv(opcode_type, 16#04#),
      2371 => to_slv(opcode_type, 16#09#),
      2372 => to_slv(opcode_type, 16#0A#),
      2373 => to_slv(opcode_type, 16#11#),
      2374 => to_slv(opcode_type, 16#07#),
      2375 => to_slv(opcode_type, 16#E2#),
      2376 => to_slv(opcode_type, 16#0A#),
      2377 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#02#),
      2402 => to_slv(opcode_type, 16#03#),
      2403 => to_slv(opcode_type, 16#05#),
      2404 => to_slv(opcode_type, 16#0D#),
      2405 => to_slv(opcode_type, 16#08#),
      2406 => to_slv(opcode_type, 16#04#),
      2407 => to_slv(opcode_type, 16#0E#),
      2408 => to_slv(opcode_type, 16#11#),
      2409 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#07#),
      2433 => to_slv(opcode_type, 16#05#),
      2434 => to_slv(opcode_type, 16#04#),
      2435 => to_slv(opcode_type, 16#01#),
      2436 => to_slv(opcode_type, 16#0F#),
      2437 => to_slv(opcode_type, 16#07#),
      2438 => to_slv(opcode_type, 16#05#),
      2439 => to_slv(opcode_type, 16#11#),
      2440 => to_slv(opcode_type, 16#0A#),
      2441 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#07#),
      2465 => to_slv(opcode_type, 16#02#),
      2466 => to_slv(opcode_type, 16#08#),
      2467 => to_slv(opcode_type, 16#08#),
      2468 => to_slv(opcode_type, 16#53#),
      2469 => to_slv(opcode_type, 16#11#),
      2470 => to_slv(opcode_type, 16#01#),
      2471 => to_slv(opcode_type, 16#10#),
      2472 => to_slv(opcode_type, 16#0D#),
      2473 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#02#),
      2497 => to_slv(opcode_type, 16#08#),
      2498 => to_slv(opcode_type, 16#07#),
      2499 => to_slv(opcode_type, 16#08#),
      2500 => to_slv(opcode_type, 16#0D#),
      2501 => to_slv(opcode_type, 16#0E#),
      2502 => to_slv(opcode_type, 16#05#),
      2503 => to_slv(opcode_type, 16#FD#),
      2504 => to_slv(opcode_type, 16#0D#),
      2505 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#04#),
      2530 => to_slv(opcode_type, 16#02#),
      2531 => to_slv(opcode_type, 16#08#),
      2532 => to_slv(opcode_type, 16#0E#),
      2533 => to_slv(opcode_type, 16#10#),
      2534 => to_slv(opcode_type, 16#07#),
      2535 => to_slv(opcode_type, 16#11#),
      2536 => to_slv(opcode_type, 16#0B#),
      2537 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#01#),
      2561 => to_slv(opcode_type, 16#02#),
      2562 => to_slv(opcode_type, 16#07#),
      2563 => to_slv(opcode_type, 16#09#),
      2564 => to_slv(opcode_type, 16#0B#),
      2565 => to_slv(opcode_type, 16#0D#),
      2566 => to_slv(opcode_type, 16#06#),
      2567 => to_slv(opcode_type, 16#0C#),
      2568 => to_slv(opcode_type, 16#0A#),
      2569 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#01#),
      2593 => to_slv(opcode_type, 16#07#),
      2594 => to_slv(opcode_type, 16#06#),
      2595 => to_slv(opcode_type, 16#03#),
      2596 => to_slv(opcode_type, 16#29#),
      2597 => to_slv(opcode_type, 16#04#),
      2598 => to_slv(opcode_type, 16#11#),
      2599 => to_slv(opcode_type, 16#03#),
      2600 => to_slv(opcode_type, 16#0F#),
      2601 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#04#),
      2625 => to_slv(opcode_type, 16#01#),
      2626 => to_slv(opcode_type, 16#06#),
      2627 => to_slv(opcode_type, 16#07#),
      2628 => to_slv(opcode_type, 16#0C#),
      2629 => to_slv(opcode_type, 16#10#),
      2630 => to_slv(opcode_type, 16#07#),
      2631 => to_slv(opcode_type, 16#11#),
      2632 => to_slv(opcode_type, 16#11#),
      2633 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#01#),
      2657 => to_slv(opcode_type, 16#07#),
      2658 => to_slv(opcode_type, 16#06#),
      2659 => to_slv(opcode_type, 16#03#),
      2660 => to_slv(opcode_type, 16#0C#),
      2661 => to_slv(opcode_type, 16#04#),
      2662 => to_slv(opcode_type, 16#0A#),
      2663 => to_slv(opcode_type, 16#01#),
      2664 => to_slv(opcode_type, 16#0C#),
      2665 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#09#),
      2689 => to_slv(opcode_type, 16#04#),
      2690 => to_slv(opcode_type, 16#02#),
      2691 => to_slv(opcode_type, 16#02#),
      2692 => to_slv(opcode_type, 16#11#),
      2693 => to_slv(opcode_type, 16#01#),
      2694 => to_slv(opcode_type, 16#05#),
      2695 => to_slv(opcode_type, 16#02#),
      2696 => to_slv(opcode_type, 16#0F#),
      2697 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#01#),
      2721 => to_slv(opcode_type, 16#08#),
      2722 => to_slv(opcode_type, 16#05#),
      2723 => to_slv(opcode_type, 16#08#),
      2724 => to_slv(opcode_type, 16#0F#),
      2725 => to_slv(opcode_type, 16#0D#),
      2726 => to_slv(opcode_type, 16#01#),
      2727 => to_slv(opcode_type, 16#05#),
      2728 => to_slv(opcode_type, 16#11#),
      2729 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#06#),
      2753 => to_slv(opcode_type, 16#05#),
      2754 => to_slv(opcode_type, 16#05#),
      2755 => to_slv(opcode_type, 16#07#),
      2756 => to_slv(opcode_type, 16#0D#),
      2757 => to_slv(opcode_type, 16#0E#),
      2758 => to_slv(opcode_type, 16#02#),
      2759 => to_slv(opcode_type, 16#04#),
      2760 => to_slv(opcode_type, 16#0A#),
      2761 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#07#),
      2785 => to_slv(opcode_type, 16#05#),
      2786 => to_slv(opcode_type, 16#03#),
      2787 => to_slv(opcode_type, 16#04#),
      2788 => to_slv(opcode_type, 16#0B#),
      2789 => to_slv(opcode_type, 16#01#),
      2790 => to_slv(opcode_type, 16#04#),
      2791 => to_slv(opcode_type, 16#02#),
      2792 => to_slv(opcode_type, 16#10#),
      2793 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#04#),
      2817 => to_slv(opcode_type, 16#08#),
      2818 => to_slv(opcode_type, 16#03#),
      2819 => to_slv(opcode_type, 16#02#),
      2820 => to_slv(opcode_type, 16#0A#),
      2821 => to_slv(opcode_type, 16#09#),
      2822 => to_slv(opcode_type, 16#01#),
      2823 => to_slv(opcode_type, 16#0E#),
      2824 => to_slv(opcode_type, 16#6D#),
      2825 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#08#),
      2849 => to_slv(opcode_type, 16#02#),
      2850 => to_slv(opcode_type, 16#02#),
      2851 => to_slv(opcode_type, 16#03#),
      2852 => to_slv(opcode_type, 16#0B#),
      2853 => to_slv(opcode_type, 16#05#),
      2854 => to_slv(opcode_type, 16#06#),
      2855 => to_slv(opcode_type, 16#0C#),
      2856 => to_slv(opcode_type, 16#0E#),
      2857 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#09#),
      2881 => to_slv(opcode_type, 16#03#),
      2882 => to_slv(opcode_type, 16#09#),
      2883 => to_slv(opcode_type, 16#03#),
      2884 => to_slv(opcode_type, 16#0D#),
      2885 => to_slv(opcode_type, 16#01#),
      2886 => to_slv(opcode_type, 16#0B#),
      2887 => to_slv(opcode_type, 16#02#),
      2888 => to_slv(opcode_type, 16#0C#),
      2889 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#03#),
      2913 => to_slv(opcode_type, 16#07#),
      2914 => to_slv(opcode_type, 16#03#),
      2915 => to_slv(opcode_type, 16#04#),
      2916 => to_slv(opcode_type, 16#0E#),
      2917 => to_slv(opcode_type, 16#09#),
      2918 => to_slv(opcode_type, 16#03#),
      2919 => to_slv(opcode_type, 16#10#),
      2920 => to_slv(opcode_type, 16#CB#),
      2921 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#08#),
      2945 => to_slv(opcode_type, 16#02#),
      2946 => to_slv(opcode_type, 16#08#),
      2947 => to_slv(opcode_type, 16#04#),
      2948 => to_slv(opcode_type, 16#0B#),
      2949 => to_slv(opcode_type, 16#02#),
      2950 => to_slv(opcode_type, 16#0A#),
      2951 => to_slv(opcode_type, 16#01#),
      2952 => to_slv(opcode_type, 16#0B#),
      2953 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#03#),
      2977 => to_slv(opcode_type, 16#02#),
      2978 => to_slv(opcode_type, 16#07#),
      2979 => to_slv(opcode_type, 16#07#),
      2980 => to_slv(opcode_type, 16#10#),
      2981 => to_slv(opcode_type, 16#0C#),
      2982 => to_slv(opcode_type, 16#06#),
      2983 => to_slv(opcode_type, 16#10#),
      2984 => to_slv(opcode_type, 16#0F#),
      2985 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#01#),
      3009 => to_slv(opcode_type, 16#07#),
      3010 => to_slv(opcode_type, 16#09#),
      3011 => to_slv(opcode_type, 16#07#),
      3012 => to_slv(opcode_type, 16#0F#),
      3013 => to_slv(opcode_type, 16#0E#),
      3014 => to_slv(opcode_type, 16#05#),
      3015 => to_slv(opcode_type, 16#11#),
      3016 => to_slv(opcode_type, 16#0B#),
      3017 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#03#),
      3041 => to_slv(opcode_type, 16#04#),
      3042 => to_slv(opcode_type, 16#09#),
      3043 => to_slv(opcode_type, 16#07#),
      3044 => to_slv(opcode_type, 16#11#),
      3045 => to_slv(opcode_type, 16#0E#),
      3046 => to_slv(opcode_type, 16#08#),
      3047 => to_slv(opcode_type, 16#0F#),
      3048 => to_slv(opcode_type, 16#0F#),
      3049 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#01#),
      3073 => to_slv(opcode_type, 16#02#),
      3074 => to_slv(opcode_type, 16#08#),
      3075 => to_slv(opcode_type, 16#08#),
      3076 => to_slv(opcode_type, 16#0C#),
      3077 => to_slv(opcode_type, 16#10#),
      3078 => to_slv(opcode_type, 16#07#),
      3079 => to_slv(opcode_type, 16#11#),
      3080 => to_slv(opcode_type, 16#11#),
      3081 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#04#),
      3105 => to_slv(opcode_type, 16#05#),
      3106 => to_slv(opcode_type, 16#09#),
      3107 => to_slv(opcode_type, 16#07#),
      3108 => to_slv(opcode_type, 16#0E#),
      3109 => to_slv(opcode_type, 16#89#),
      3110 => to_slv(opcode_type, 16#08#),
      3111 => to_slv(opcode_type, 16#0B#),
      3112 => to_slv(opcode_type, 16#0B#),
      3113 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#05#),
      3137 => to_slv(opcode_type, 16#09#),
      3138 => to_slv(opcode_type, 16#02#),
      3139 => to_slv(opcode_type, 16#07#),
      3140 => to_slv(opcode_type, 16#0D#),
      3141 => to_slv(opcode_type, 16#0B#),
      3142 => to_slv(opcode_type, 16#05#),
      3143 => to_slv(opcode_type, 16#03#),
      3144 => to_slv(opcode_type, 16#0C#),
      3145 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#07#),
      3169 => to_slv(opcode_type, 16#07#),
      3170 => to_slv(opcode_type, 16#04#),
      3171 => to_slv(opcode_type, 16#01#),
      3172 => to_slv(opcode_type, 16#0F#),
      3173 => to_slv(opcode_type, 16#08#),
      3174 => to_slv(opcode_type, 16#C2#),
      3175 => to_slv(opcode_type, 16#0D#),
      3176 => to_slv(opcode_type, 16#10#),
      3177 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#03#),
      3201 => to_slv(opcode_type, 16#05#),
      3202 => to_slv(opcode_type, 16#09#),
      3203 => to_slv(opcode_type, 16#09#),
      3204 => to_slv(opcode_type, 16#0C#),
      3205 => to_slv(opcode_type, 16#5E#),
      3206 => to_slv(opcode_type, 16#07#),
      3207 => to_slv(opcode_type, 16#0B#),
      3208 => to_slv(opcode_type, 16#0A#),
      3209 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#04#),
      3233 => to_slv(opcode_type, 16#09#),
      3234 => to_slv(opcode_type, 16#02#),
      3235 => to_slv(opcode_type, 16#05#),
      3236 => to_slv(opcode_type, 16#0A#),
      3237 => to_slv(opcode_type, 16#07#),
      3238 => to_slv(opcode_type, 16#02#),
      3239 => to_slv(opcode_type, 16#0C#),
      3240 => to_slv(opcode_type, 16#45#),
      3241 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#01#),
      3265 => to_slv(opcode_type, 16#04#),
      3266 => to_slv(opcode_type, 16#07#),
      3267 => to_slv(opcode_type, 16#06#),
      3268 => to_slv(opcode_type, 16#0D#),
      3269 => to_slv(opcode_type, 16#A5#),
      3270 => to_slv(opcode_type, 16#07#),
      3271 => to_slv(opcode_type, 16#0D#),
      3272 => to_slv(opcode_type, 16#0D#),
      3273 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#02#),
      3297 => to_slv(opcode_type, 16#07#),
      3298 => to_slv(opcode_type, 16#03#),
      3299 => to_slv(opcode_type, 16#06#),
      3300 => to_slv(opcode_type, 16#0D#),
      3301 => to_slv(opcode_type, 16#0D#),
      3302 => to_slv(opcode_type, 16#07#),
      3303 => to_slv(opcode_type, 16#0D#),
      3304 => to_slv(opcode_type, 16#10#),
      3305 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#08#),
      3329 => to_slv(opcode_type, 16#07#),
      3330 => to_slv(opcode_type, 16#07#),
      3331 => to_slv(opcode_type, 16#05#),
      3332 => to_slv(opcode_type, 16#0B#),
      3333 => to_slv(opcode_type, 16#01#),
      3334 => to_slv(opcode_type, 16#0B#),
      3335 => to_slv(opcode_type, 16#0E#),
      3336 => to_slv(opcode_type, 16#11#),
      3337 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#01#),
      3361 => to_slv(opcode_type, 16#04#),
      3362 => to_slv(opcode_type, 16#06#),
      3363 => to_slv(opcode_type, 16#08#),
      3364 => to_slv(opcode_type, 16#0E#),
      3365 => to_slv(opcode_type, 16#0F#),
      3366 => to_slv(opcode_type, 16#08#),
      3367 => to_slv(opcode_type, 16#0F#),
      3368 => to_slv(opcode_type, 16#10#),
      3369 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#03#),
      3393 => to_slv(opcode_type, 16#06#),
      3394 => to_slv(opcode_type, 16#08#),
      3395 => to_slv(opcode_type, 16#02#),
      3396 => to_slv(opcode_type, 16#F0#),
      3397 => to_slv(opcode_type, 16#06#),
      3398 => to_slv(opcode_type, 16#10#),
      3399 => to_slv(opcode_type, 16#0C#),
      3400 => to_slv(opcode_type, 16#0F#),
      3401 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#02#),
      3426 => to_slv(opcode_type, 16#03#),
      3427 => to_slv(opcode_type, 16#06#),
      3428 => to_slv(opcode_type, 16#0C#),
      3429 => to_slv(opcode_type, 16#0F#),
      3430 => to_slv(opcode_type, 16#02#),
      3431 => to_slv(opcode_type, 16#04#),
      3432 => to_slv(opcode_type, 16#0D#),
      3433 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#04#),
      3457 => to_slv(opcode_type, 16#01#),
      3458 => to_slv(opcode_type, 16#09#),
      3459 => to_slv(opcode_type, 16#09#),
      3460 => to_slv(opcode_type, 16#0A#),
      3461 => to_slv(opcode_type, 16#11#),
      3462 => to_slv(opcode_type, 16#06#),
      3463 => to_slv(opcode_type, 16#11#),
      3464 => to_slv(opcode_type, 16#0B#),
      3465 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#03#),
      3489 => to_slv(opcode_type, 16#09#),
      3490 => to_slv(opcode_type, 16#04#),
      3491 => to_slv(opcode_type, 16#09#),
      3492 => to_slv(opcode_type, 16#0C#),
      3493 => to_slv(opcode_type, 16#0B#),
      3494 => to_slv(opcode_type, 16#06#),
      3495 => to_slv(opcode_type, 16#20#),
      3496 => to_slv(opcode_type, 16#0F#),
      3497 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#08#),
      3521 => to_slv(opcode_type, 16#08#),
      3522 => to_slv(opcode_type, 16#08#),
      3523 => to_slv(opcode_type, 16#04#),
      3524 => to_slv(opcode_type, 16#0B#),
      3525 => to_slv(opcode_type, 16#04#),
      3526 => to_slv(opcode_type, 16#50#),
      3527 => to_slv(opcode_type, 16#10#),
      3528 => to_slv(opcode_type, 16#0F#),
      3529 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#08#),
      3553 => to_slv(opcode_type, 16#04#),
      3554 => to_slv(opcode_type, 16#03#),
      3555 => to_slv(opcode_type, 16#06#),
      3556 => to_slv(opcode_type, 16#0F#),
      3557 => to_slv(opcode_type, 16#0F#),
      3558 => to_slv(opcode_type, 16#02#),
      3559 => to_slv(opcode_type, 16#01#),
      3560 => to_slv(opcode_type, 16#0E#),
      3561 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#07#),
      3585 => to_slv(opcode_type, 16#03#),
      3586 => to_slv(opcode_type, 16#03#),
      3587 => to_slv(opcode_type, 16#07#),
      3588 => to_slv(opcode_type, 16#10#),
      3589 => to_slv(opcode_type, 16#0B#),
      3590 => to_slv(opcode_type, 16#02#),
      3591 => to_slv(opcode_type, 16#05#),
      3592 => to_slv(opcode_type, 16#0F#),
      3593 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#04#),
      3617 => to_slv(opcode_type, 16#09#),
      3618 => to_slv(opcode_type, 16#02#),
      3619 => to_slv(opcode_type, 16#06#),
      3620 => to_slv(opcode_type, 16#0C#),
      3621 => to_slv(opcode_type, 16#0F#),
      3622 => to_slv(opcode_type, 16#05#),
      3623 => to_slv(opcode_type, 16#03#),
      3624 => to_slv(opcode_type, 16#AB#),
      3625 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#01#),
      3649 => to_slv(opcode_type, 16#05#),
      3650 => to_slv(opcode_type, 16#07#),
      3651 => to_slv(opcode_type, 16#09#),
      3652 => to_slv(opcode_type, 16#0B#),
      3653 => to_slv(opcode_type, 16#11#),
      3654 => to_slv(opcode_type, 16#09#),
      3655 => to_slv(opcode_type, 16#11#),
      3656 => to_slv(opcode_type, 16#0B#),
      3657 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#01#),
      3681 => to_slv(opcode_type, 16#07#),
      3682 => to_slv(opcode_type, 16#08#),
      3683 => to_slv(opcode_type, 16#06#),
      3684 => to_slv(opcode_type, 16#0C#),
      3685 => to_slv(opcode_type, 16#0A#),
      3686 => to_slv(opcode_type, 16#03#),
      3687 => to_slv(opcode_type, 16#0B#),
      3688 => to_slv(opcode_type, 16#0C#),
      3689 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#01#),
      3713 => to_slv(opcode_type, 16#02#),
      3714 => to_slv(opcode_type, 16#09#),
      3715 => to_slv(opcode_type, 16#08#),
      3716 => to_slv(opcode_type, 16#0D#),
      3717 => to_slv(opcode_type, 16#0F#),
      3718 => to_slv(opcode_type, 16#06#),
      3719 => to_slv(opcode_type, 16#10#),
      3720 => to_slv(opcode_type, 16#0E#),
      3721 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#01#),
      3745 => to_slv(opcode_type, 16#02#),
      3746 => to_slv(opcode_type, 16#06#),
      3747 => to_slv(opcode_type, 16#06#),
      3748 => to_slv(opcode_type, 16#10#),
      3749 => to_slv(opcode_type, 16#3E#),
      3750 => to_slv(opcode_type, 16#06#),
      3751 => to_slv(opcode_type, 16#0F#),
      3752 => to_slv(opcode_type, 16#11#),
      3753 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#04#),
      3777 => to_slv(opcode_type, 16#04#),
      3778 => to_slv(opcode_type, 16#08#),
      3779 => to_slv(opcode_type, 16#08#),
      3780 => to_slv(opcode_type, 16#3A#),
      3781 => to_slv(opcode_type, 16#10#),
      3782 => to_slv(opcode_type, 16#06#),
      3783 => to_slv(opcode_type, 16#BD#),
      3784 => to_slv(opcode_type, 16#0E#),
      3785 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#05#),
      3809 => to_slv(opcode_type, 16#06#),
      3810 => to_slv(opcode_type, 16#03#),
      3811 => to_slv(opcode_type, 16#02#),
      3812 => to_slv(opcode_type, 16#0D#),
      3813 => to_slv(opcode_type, 16#02#),
      3814 => to_slv(opcode_type, 16#07#),
      3815 => to_slv(opcode_type, 16#FF#),
      3816 => to_slv(opcode_type, 16#0A#),
      3817 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#08#),
      3841 => to_slv(opcode_type, 16#08#),
      3842 => to_slv(opcode_type, 16#01#),
      3843 => to_slv(opcode_type, 16#09#),
      3844 => to_slv(opcode_type, 16#0B#),
      3845 => to_slv(opcode_type, 16#0B#),
      3846 => to_slv(opcode_type, 16#02#),
      3847 => to_slv(opcode_type, 16#0B#),
      3848 => to_slv(opcode_type, 16#0B#),
      3849 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#08#),
      3873 => to_slv(opcode_type, 16#04#),
      3874 => to_slv(opcode_type, 16#01#),
      3875 => to_slv(opcode_type, 16#08#),
      3876 => to_slv(opcode_type, 16#0E#),
      3877 => to_slv(opcode_type, 16#0B#),
      3878 => to_slv(opcode_type, 16#08#),
      3879 => to_slv(opcode_type, 16#0E#),
      3880 => to_slv(opcode_type, 16#0C#),
      3881 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#08#),
      3905 => to_slv(opcode_type, 16#07#),
      3906 => to_slv(opcode_type, 16#03#),
      3907 => to_slv(opcode_type, 16#07#),
      3908 => to_slv(opcode_type, 16#13#),
      3909 => to_slv(opcode_type, 16#0A#),
      3910 => to_slv(opcode_type, 16#01#),
      3911 => to_slv(opcode_type, 16#0B#),
      3912 => to_slv(opcode_type, 16#11#),
      3913 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#04#),
      3937 => to_slv(opcode_type, 16#05#),
      3938 => to_slv(opcode_type, 16#06#),
      3939 => to_slv(opcode_type, 16#08#),
      3940 => to_slv(opcode_type, 16#0A#),
      3941 => to_slv(opcode_type, 16#0A#),
      3942 => to_slv(opcode_type, 16#07#),
      3943 => to_slv(opcode_type, 16#0F#),
      3944 => to_slv(opcode_type, 16#10#),
      3945 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#04#),
      3969 => to_slv(opcode_type, 16#02#),
      3970 => to_slv(opcode_type, 16#09#),
      3971 => to_slv(opcode_type, 16#08#),
      3972 => to_slv(opcode_type, 16#0F#),
      3973 => to_slv(opcode_type, 16#0D#),
      3974 => to_slv(opcode_type, 16#08#),
      3975 => to_slv(opcode_type, 16#0E#),
      3976 => to_slv(opcode_type, 16#0A#),
      3977 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#02#),
      4001 => to_slv(opcode_type, 16#07#),
      4002 => to_slv(opcode_type, 16#05#),
      4003 => to_slv(opcode_type, 16#03#),
      4004 => to_slv(opcode_type, 16#10#),
      4005 => to_slv(opcode_type, 16#07#),
      4006 => to_slv(opcode_type, 16#01#),
      4007 => to_slv(opcode_type, 16#0F#),
      4008 => to_slv(opcode_type, 16#6F#),
      4009 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#03#),
      4033 => to_slv(opcode_type, 16#08#),
      4034 => to_slv(opcode_type, 16#04#),
      4035 => to_slv(opcode_type, 16#06#),
      4036 => to_slv(opcode_type, 16#0F#),
      4037 => to_slv(opcode_type, 16#0A#),
      4038 => to_slv(opcode_type, 16#02#),
      4039 => to_slv(opcode_type, 16#01#),
      4040 => to_slv(opcode_type, 16#0B#),
      4041 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#05#),
      4065 => to_slv(opcode_type, 16#06#),
      4066 => to_slv(opcode_type, 16#06#),
      4067 => to_slv(opcode_type, 16#01#),
      4068 => to_slv(opcode_type, 16#11#),
      4069 => to_slv(opcode_type, 16#01#),
      4070 => to_slv(opcode_type, 16#0A#),
      4071 => to_slv(opcode_type, 16#04#),
      4072 => to_slv(opcode_type, 16#0C#),
      4073 to 4095 => (others => '0')
  ),

    -- Bin `10`...
    9 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#04#),
      1 => to_slv(opcode_type, 16#09#),
      2 => to_slv(opcode_type, 16#07#),
      3 => to_slv(opcode_type, 16#06#),
      4 => to_slv(opcode_type, 16#0F#),
      5 => to_slv(opcode_type, 16#0C#),
      6 => to_slv(opcode_type, 16#05#),
      7 => to_slv(opcode_type, 16#0D#),
      8 => to_slv(opcode_type, 16#03#),
      9 => to_slv(opcode_type, 16#0D#),
      10 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#01#),
      33 => to_slv(opcode_type, 16#09#),
      34 => to_slv(opcode_type, 16#05#),
      35 => to_slv(opcode_type, 16#05#),
      36 => to_slv(opcode_type, 16#0B#),
      37 => to_slv(opcode_type, 16#07#),
      38 => to_slv(opcode_type, 16#05#),
      39 => to_slv(opcode_type, 16#11#),
      40 => to_slv(opcode_type, 16#01#),
      41 => to_slv(opcode_type, 16#0F#),
      42 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#08#),
      65 => to_slv(opcode_type, 16#02#),
      66 => to_slv(opcode_type, 16#07#),
      67 => to_slv(opcode_type, 16#02#),
      68 => to_slv(opcode_type, 16#0E#),
      69 => to_slv(opcode_type, 16#07#),
      70 => to_slv(opcode_type, 16#10#),
      71 => to_slv(opcode_type, 16#0C#),
      72 => to_slv(opcode_type, 16#05#),
      73 => to_slv(opcode_type, 16#11#),
      74 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#07#),
      97 => to_slv(opcode_type, 16#01#),
      98 => to_slv(opcode_type, 16#04#),
      99 => to_slv(opcode_type, 16#03#),
      100 => to_slv(opcode_type, 16#0C#),
      101 => to_slv(opcode_type, 16#05#),
      102 => to_slv(opcode_type, 16#07#),
      103 => to_slv(opcode_type, 16#03#),
      104 => to_slv(opcode_type, 16#0C#),
      105 => to_slv(opcode_type, 16#0D#),
      106 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#03#),
      129 => to_slv(opcode_type, 16#09#),
      130 => to_slv(opcode_type, 16#04#),
      131 => to_slv(opcode_type, 16#09#),
      132 => to_slv(opcode_type, 16#0A#),
      133 => to_slv(opcode_type, 16#0E#),
      134 => to_slv(opcode_type, 16#09#),
      135 => to_slv(opcode_type, 16#04#),
      136 => to_slv(opcode_type, 16#B6#),
      137 => to_slv(opcode_type, 16#CD#),
      138 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#06#),
      161 => to_slv(opcode_type, 16#06#),
      162 => to_slv(opcode_type, 16#08#),
      163 => to_slv(opcode_type, 16#05#),
      164 => to_slv(opcode_type, 16#0B#),
      165 => to_slv(opcode_type, 16#04#),
      166 => to_slv(opcode_type, 16#C8#),
      167 => to_slv(opcode_type, 16#01#),
      168 => to_slv(opcode_type, 16#0B#),
      169 => to_slv(opcode_type, 16#0E#),
      170 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#03#),
      193 => to_slv(opcode_type, 16#07#),
      194 => to_slv(opcode_type, 16#03#),
      195 => to_slv(opcode_type, 16#05#),
      196 => to_slv(opcode_type, 16#0C#),
      197 => to_slv(opcode_type, 16#09#),
      198 => to_slv(opcode_type, 16#03#),
      199 => to_slv(opcode_type, 16#0A#),
      200 => to_slv(opcode_type, 16#04#),
      201 => to_slv(opcode_type, 16#0F#),
      202 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#02#),
      225 => to_slv(opcode_type, 16#08#),
      226 => to_slv(opcode_type, 16#07#),
      227 => to_slv(opcode_type, 16#03#),
      228 => to_slv(opcode_type, 16#16#),
      229 => to_slv(opcode_type, 16#06#),
      230 => to_slv(opcode_type, 16#0E#),
      231 => to_slv(opcode_type, 16#8D#),
      232 => to_slv(opcode_type, 16#05#),
      233 => to_slv(opcode_type, 16#0A#),
      234 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#01#),
      257 => to_slv(opcode_type, 16#06#),
      258 => to_slv(opcode_type, 16#09#),
      259 => to_slv(opcode_type, 16#05#),
      260 => to_slv(opcode_type, 16#10#),
      261 => to_slv(opcode_type, 16#02#),
      262 => to_slv(opcode_type, 16#10#),
      263 => to_slv(opcode_type, 16#05#),
      264 => to_slv(opcode_type, 16#02#),
      265 => to_slv(opcode_type, 16#0E#),
      266 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#04#),
      289 => to_slv(opcode_type, 16#06#),
      290 => to_slv(opcode_type, 16#06#),
      291 => to_slv(opcode_type, 16#09#),
      292 => to_slv(opcode_type, 16#0A#),
      293 => to_slv(opcode_type, 16#10#),
      294 => to_slv(opcode_type, 16#07#),
      295 => to_slv(opcode_type, 16#26#),
      296 => to_slv(opcode_type, 16#0A#),
      297 => to_slv(opcode_type, 16#11#),
      298 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#06#),
      321 => to_slv(opcode_type, 16#03#),
      322 => to_slv(opcode_type, 16#01#),
      323 => to_slv(opcode_type, 16#04#),
      324 => to_slv(opcode_type, 16#0D#),
      325 => to_slv(opcode_type, 16#07#),
      326 => to_slv(opcode_type, 16#02#),
      327 => to_slv(opcode_type, 16#04#),
      328 => to_slv(opcode_type, 16#0A#),
      329 => to_slv(opcode_type, 16#0E#),
      330 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#07#),
      353 => to_slv(opcode_type, 16#08#),
      354 => to_slv(opcode_type, 16#01#),
      355 => to_slv(opcode_type, 16#04#),
      356 => to_slv(opcode_type, 16#0F#),
      357 => to_slv(opcode_type, 16#02#),
      358 => to_slv(opcode_type, 16#05#),
      359 => to_slv(opcode_type, 16#0D#),
      360 => to_slv(opcode_type, 16#03#),
      361 => to_slv(opcode_type, 16#0C#),
      362 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#01#),
      385 => to_slv(opcode_type, 16#06#),
      386 => to_slv(opcode_type, 16#07#),
      387 => to_slv(opcode_type, 16#09#),
      388 => to_slv(opcode_type, 16#0C#),
      389 => to_slv(opcode_type, 16#0F#),
      390 => to_slv(opcode_type, 16#02#),
      391 => to_slv(opcode_type, 16#0D#),
      392 => to_slv(opcode_type, 16#05#),
      393 => to_slv(opcode_type, 16#0A#),
      394 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#01#),
      417 => to_slv(opcode_type, 16#06#),
      418 => to_slv(opcode_type, 16#08#),
      419 => to_slv(opcode_type, 16#08#),
      420 => to_slv(opcode_type, 16#0D#),
      421 => to_slv(opcode_type, 16#0E#),
      422 => to_slv(opcode_type, 16#06#),
      423 => to_slv(opcode_type, 16#0E#),
      424 => to_slv(opcode_type, 16#0C#),
      425 => to_slv(opcode_type, 16#10#),
      426 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#03#),
      449 => to_slv(opcode_type, 16#06#),
      450 => to_slv(opcode_type, 16#01#),
      451 => to_slv(opcode_type, 16#03#),
      452 => to_slv(opcode_type, 16#0D#),
      453 => to_slv(opcode_type, 16#08#),
      454 => to_slv(opcode_type, 16#02#),
      455 => to_slv(opcode_type, 16#0D#),
      456 => to_slv(opcode_type, 16#05#),
      457 => to_slv(opcode_type, 16#0E#),
      458 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#02#),
      481 => to_slv(opcode_type, 16#06#),
      482 => to_slv(opcode_type, 16#01#),
      483 => to_slv(opcode_type, 16#04#),
      484 => to_slv(opcode_type, 16#0E#),
      485 => to_slv(opcode_type, 16#06#),
      486 => to_slv(opcode_type, 16#02#),
      487 => to_slv(opcode_type, 16#0B#),
      488 => to_slv(opcode_type, 16#01#),
      489 => to_slv(opcode_type, 16#0B#),
      490 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#09#),
      514 => to_slv(opcode_type, 16#08#),
      515 => to_slv(opcode_type, 16#08#),
      516 => to_slv(opcode_type, 16#0B#),
      517 => to_slv(opcode_type, 16#10#),
      518 => to_slv(opcode_type, 16#05#),
      519 => to_slv(opcode_type, 16#10#),
      520 => to_slv(opcode_type, 16#0D#),
      521 => to_slv(opcode_type, 16#0D#),
      522 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#05#),
      545 => to_slv(opcode_type, 16#07#),
      546 => to_slv(opcode_type, 16#03#),
      547 => to_slv(opcode_type, 16#08#),
      548 => to_slv(opcode_type, 16#10#),
      549 => to_slv(opcode_type, 16#0A#),
      550 => to_slv(opcode_type, 16#09#),
      551 => to_slv(opcode_type, 16#02#),
      552 => to_slv(opcode_type, 16#0E#),
      553 => to_slv(opcode_type, 16#0A#),
      554 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#04#),
      577 => to_slv(opcode_type, 16#07#),
      578 => to_slv(opcode_type, 16#05#),
      579 => to_slv(opcode_type, 16#03#),
      580 => to_slv(opcode_type, 16#0B#),
      581 => to_slv(opcode_type, 16#07#),
      582 => to_slv(opcode_type, 16#03#),
      583 => to_slv(opcode_type, 16#0A#),
      584 => to_slv(opcode_type, 16#04#),
      585 => to_slv(opcode_type, 16#11#),
      586 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#04#),
      609 => to_slv(opcode_type, 16#06#),
      610 => to_slv(opcode_type, 16#02#),
      611 => to_slv(opcode_type, 16#02#),
      612 => to_slv(opcode_type, 16#10#),
      613 => to_slv(opcode_type, 16#06#),
      614 => to_slv(opcode_type, 16#07#),
      615 => to_slv(opcode_type, 16#11#),
      616 => to_slv(opcode_type, 16#10#),
      617 => to_slv(opcode_type, 16#0B#),
      618 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#05#),
      641 => to_slv(opcode_type, 16#08#),
      642 => to_slv(opcode_type, 16#05#),
      643 => to_slv(opcode_type, 16#04#),
      644 => to_slv(opcode_type, 16#0D#),
      645 => to_slv(opcode_type, 16#09#),
      646 => to_slv(opcode_type, 16#08#),
      647 => to_slv(opcode_type, 16#0F#),
      648 => to_slv(opcode_type, 16#0A#),
      649 => to_slv(opcode_type, 16#0B#),
      650 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#07#),
      673 => to_slv(opcode_type, 16#07#),
      674 => to_slv(opcode_type, 16#05#),
      675 => to_slv(opcode_type, 16#07#),
      676 => to_slv(opcode_type, 16#10#),
      677 => to_slv(opcode_type, 16#0A#),
      678 => to_slv(opcode_type, 16#05#),
      679 => to_slv(opcode_type, 16#03#),
      680 => to_slv(opcode_type, 16#C9#),
      681 => to_slv(opcode_type, 16#10#),
      682 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#02#),
      705 => to_slv(opcode_type, 16#09#),
      706 => to_slv(opcode_type, 16#03#),
      707 => to_slv(opcode_type, 16#08#),
      708 => to_slv(opcode_type, 16#10#),
      709 => to_slv(opcode_type, 16#78#),
      710 => to_slv(opcode_type, 16#06#),
      711 => to_slv(opcode_type, 16#02#),
      712 => to_slv(opcode_type, 16#0E#),
      713 => to_slv(opcode_type, 16#0C#),
      714 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#02#),
      737 => to_slv(opcode_type, 16#06#),
      738 => to_slv(opcode_type, 16#08#),
      739 => to_slv(opcode_type, 16#03#),
      740 => to_slv(opcode_type, 16#0F#),
      741 => to_slv(opcode_type, 16#07#),
      742 => to_slv(opcode_type, 16#0A#),
      743 => to_slv(opcode_type, 16#72#),
      744 => to_slv(opcode_type, 16#05#),
      745 => to_slv(opcode_type, 16#10#),
      746 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#02#),
      769 => to_slv(opcode_type, 16#09#),
      770 => to_slv(opcode_type, 16#09#),
      771 => to_slv(opcode_type, 16#01#),
      772 => to_slv(opcode_type, 16#0E#),
      773 => to_slv(opcode_type, 16#03#),
      774 => to_slv(opcode_type, 16#0A#),
      775 => to_slv(opcode_type, 16#02#),
      776 => to_slv(opcode_type, 16#01#),
      777 => to_slv(opcode_type, 16#0F#),
      778 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#05#),
      801 => to_slv(opcode_type, 16#08#),
      802 => to_slv(opcode_type, 16#05#),
      803 => to_slv(opcode_type, 16#04#),
      804 => to_slv(opcode_type, 16#0B#),
      805 => to_slv(opcode_type, 16#07#),
      806 => to_slv(opcode_type, 16#08#),
      807 => to_slv(opcode_type, 16#0D#),
      808 => to_slv(opcode_type, 16#11#),
      809 => to_slv(opcode_type, 16#11#),
      810 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#07#),
      833 => to_slv(opcode_type, 16#05#),
      834 => to_slv(opcode_type, 16#08#),
      835 => to_slv(opcode_type, 16#03#),
      836 => to_slv(opcode_type, 16#0F#),
      837 => to_slv(opcode_type, 16#03#),
      838 => to_slv(opcode_type, 16#0C#),
      839 => to_slv(opcode_type, 16#02#),
      840 => to_slv(opcode_type, 16#05#),
      841 => to_slv(opcode_type, 16#0F#),
      842 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#06#),
      865 => to_slv(opcode_type, 16#08#),
      866 => to_slv(opcode_type, 16#09#),
      867 => to_slv(opcode_type, 16#06#),
      868 => to_slv(opcode_type, 16#0F#),
      869 => to_slv(opcode_type, 16#0D#),
      870 => to_slv(opcode_type, 16#01#),
      871 => to_slv(opcode_type, 16#40#),
      872 => to_slv(opcode_type, 16#0F#),
      873 => to_slv(opcode_type, 16#0C#),
      874 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#04#),
      897 => to_slv(opcode_type, 16#09#),
      898 => to_slv(opcode_type, 16#01#),
      899 => to_slv(opcode_type, 16#07#),
      900 => to_slv(opcode_type, 16#0D#),
      901 => to_slv(opcode_type, 16#0E#),
      902 => to_slv(opcode_type, 16#08#),
      903 => to_slv(opcode_type, 16#04#),
      904 => to_slv(opcode_type, 16#0B#),
      905 => to_slv(opcode_type, 16#0D#),
      906 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#03#),
      929 => to_slv(opcode_type, 16#07#),
      930 => to_slv(opcode_type, 16#05#),
      931 => to_slv(opcode_type, 16#03#),
      932 => to_slv(opcode_type, 16#7C#),
      933 => to_slv(opcode_type, 16#09#),
      934 => to_slv(opcode_type, 16#03#),
      935 => to_slv(opcode_type, 16#0E#),
      936 => to_slv(opcode_type, 16#05#),
      937 => to_slv(opcode_type, 16#0F#),
      938 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#01#),
      961 => to_slv(opcode_type, 16#07#),
      962 => to_slv(opcode_type, 16#04#),
      963 => to_slv(opcode_type, 16#05#),
      964 => to_slv(opcode_type, 16#0C#),
      965 => to_slv(opcode_type, 16#06#),
      966 => to_slv(opcode_type, 16#03#),
      967 => to_slv(opcode_type, 16#0E#),
      968 => to_slv(opcode_type, 16#02#),
      969 => to_slv(opcode_type, 16#10#),
      970 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#02#),
      993 => to_slv(opcode_type, 16#09#),
      994 => to_slv(opcode_type, 16#08#),
      995 => to_slv(opcode_type, 16#01#),
      996 => to_slv(opcode_type, 16#0D#),
      997 => to_slv(opcode_type, 16#09#),
      998 => to_slv(opcode_type, 16#11#),
      999 => to_slv(opcode_type, 16#0C#),
      1000 => to_slv(opcode_type, 16#03#),
      1001 => to_slv(opcode_type, 16#10#),
      1002 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#01#),
      1025 => to_slv(opcode_type, 16#08#),
      1026 => to_slv(opcode_type, 16#05#),
      1027 => to_slv(opcode_type, 16#01#),
      1028 => to_slv(opcode_type, 16#10#),
      1029 => to_slv(opcode_type, 16#06#),
      1030 => to_slv(opcode_type, 16#08#),
      1031 => to_slv(opcode_type, 16#10#),
      1032 => to_slv(opcode_type, 16#11#),
      1033 => to_slv(opcode_type, 16#10#),
      1034 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#08#),
      1057 => to_slv(opcode_type, 16#06#),
      1058 => to_slv(opcode_type, 16#03#),
      1059 => to_slv(opcode_type, 16#07#),
      1060 => to_slv(opcode_type, 16#0C#),
      1061 => to_slv(opcode_type, 16#0F#),
      1062 => to_slv(opcode_type, 16#09#),
      1063 => to_slv(opcode_type, 16#34#),
      1064 => to_slv(opcode_type, 16#10#),
      1065 => to_slv(opcode_type, 16#0A#),
      1066 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#01#),
      1089 => to_slv(opcode_type, 16#08#),
      1090 => to_slv(opcode_type, 16#06#),
      1091 => to_slv(opcode_type, 16#05#),
      1092 => to_slv(opcode_type, 16#0C#),
      1093 => to_slv(opcode_type, 16#04#),
      1094 => to_slv(opcode_type, 16#0A#),
      1095 => to_slv(opcode_type, 16#08#),
      1096 => to_slv(opcode_type, 16#90#),
      1097 => to_slv(opcode_type, 16#0E#),
      1098 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#07#),
      1121 => to_slv(opcode_type, 16#04#),
      1122 => to_slv(opcode_type, 16#09#),
      1123 => to_slv(opcode_type, 16#03#),
      1124 => to_slv(opcode_type, 16#0F#),
      1125 => to_slv(opcode_type, 16#09#),
      1126 => to_slv(opcode_type, 16#0C#),
      1127 => to_slv(opcode_type, 16#10#),
      1128 => to_slv(opcode_type, 16#03#),
      1129 => to_slv(opcode_type, 16#11#),
      1130 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#05#),
      1153 => to_slv(opcode_type, 16#06#),
      1154 => to_slv(opcode_type, 16#06#),
      1155 => to_slv(opcode_type, 16#08#),
      1156 => to_slv(opcode_type, 16#3C#),
      1157 => to_slv(opcode_type, 16#11#),
      1158 => to_slv(opcode_type, 16#02#),
      1159 => to_slv(opcode_type, 16#0C#),
      1160 => to_slv(opcode_type, 16#04#),
      1161 => to_slv(opcode_type, 16#11#),
      1162 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#04#),
      1185 => to_slv(opcode_type, 16#06#),
      1186 => to_slv(opcode_type, 16#07#),
      1187 => to_slv(opcode_type, 16#06#),
      1188 => to_slv(opcode_type, 16#0F#),
      1189 => to_slv(opcode_type, 16#0F#),
      1190 => to_slv(opcode_type, 16#01#),
      1191 => to_slv(opcode_type, 16#0F#),
      1192 => to_slv(opcode_type, 16#02#),
      1193 => to_slv(opcode_type, 16#0F#),
      1194 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#01#),
      1217 => to_slv(opcode_type, 16#07#),
      1218 => to_slv(opcode_type, 16#04#),
      1219 => to_slv(opcode_type, 16#08#),
      1220 => to_slv(opcode_type, 16#10#),
      1221 => to_slv(opcode_type, 16#0C#),
      1222 => to_slv(opcode_type, 16#02#),
      1223 => to_slv(opcode_type, 16#07#),
      1224 => to_slv(opcode_type, 16#10#),
      1225 => to_slv(opcode_type, 16#0A#),
      1226 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#09#),
      1249 => to_slv(opcode_type, 16#07#),
      1250 => to_slv(opcode_type, 16#06#),
      1251 => to_slv(opcode_type, 16#04#),
      1252 => to_slv(opcode_type, 16#0F#),
      1253 => to_slv(opcode_type, 16#04#),
      1254 => to_slv(opcode_type, 16#96#),
      1255 => to_slv(opcode_type, 16#01#),
      1256 => to_slv(opcode_type, 16#10#),
      1257 => to_slv(opcode_type, 16#0E#),
      1258 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#03#),
      1282 => to_slv(opcode_type, 16#07#),
      1283 => to_slv(opcode_type, 16#08#),
      1284 => to_slv(opcode_type, 16#0D#),
      1285 => to_slv(opcode_type, 16#0A#),
      1286 => to_slv(opcode_type, 16#09#),
      1287 => to_slv(opcode_type, 16#0D#),
      1288 => to_slv(opcode_type, 16#0C#),
      1289 => to_slv(opcode_type, 16#0D#),
      1290 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#03#),
      1313 => to_slv(opcode_type, 16#09#),
      1314 => to_slv(opcode_type, 16#02#),
      1315 => to_slv(opcode_type, 16#05#),
      1316 => to_slv(opcode_type, 16#10#),
      1317 => to_slv(opcode_type, 16#07#),
      1318 => to_slv(opcode_type, 16#06#),
      1319 => to_slv(opcode_type, 16#0D#),
      1320 => to_slv(opcode_type, 16#10#),
      1321 => to_slv(opcode_type, 16#10#),
      1322 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#02#),
      1345 => to_slv(opcode_type, 16#07#),
      1346 => to_slv(opcode_type, 16#05#),
      1347 => to_slv(opcode_type, 16#03#),
      1348 => to_slv(opcode_type, 16#10#),
      1349 => to_slv(opcode_type, 16#06#),
      1350 => to_slv(opcode_type, 16#05#),
      1351 => to_slv(opcode_type, 16#0B#),
      1352 => to_slv(opcode_type, 16#04#),
      1353 => to_slv(opcode_type, 16#11#),
      1354 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#09#),
      1377 => to_slv(opcode_type, 16#01#),
      1378 => to_slv(opcode_type, 16#01#),
      1379 => to_slv(opcode_type, 16#05#),
      1380 => to_slv(opcode_type, 16#0B#),
      1381 => to_slv(opcode_type, 16#05#),
      1382 => to_slv(opcode_type, 16#05#),
      1383 => to_slv(opcode_type, 16#07#),
      1384 => to_slv(opcode_type, 16#0A#),
      1385 => to_slv(opcode_type, 16#0A#),
      1386 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#09#),
      1409 => to_slv(opcode_type, 16#06#),
      1410 => to_slv(opcode_type, 16#02#),
      1411 => to_slv(opcode_type, 16#02#),
      1412 => to_slv(opcode_type, 16#0F#),
      1413 => to_slv(opcode_type, 16#02#),
      1414 => to_slv(opcode_type, 16#03#),
      1415 => to_slv(opcode_type, 16#11#),
      1416 => to_slv(opcode_type, 16#02#),
      1417 => to_slv(opcode_type, 16#10#),
      1418 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#08#),
      1441 => to_slv(opcode_type, 16#02#),
      1442 => to_slv(opcode_type, 16#07#),
      1443 => to_slv(opcode_type, 16#03#),
      1444 => to_slv(opcode_type, 16#0D#),
      1445 => to_slv(opcode_type, 16#06#),
      1446 => to_slv(opcode_type, 16#11#),
      1447 => to_slv(opcode_type, 16#0C#),
      1448 => to_slv(opcode_type, 16#01#),
      1449 => to_slv(opcode_type, 16#11#),
      1450 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#09#),
      1473 => to_slv(opcode_type, 16#08#),
      1474 => to_slv(opcode_type, 16#06#),
      1475 => to_slv(opcode_type, 16#06#),
      1476 => to_slv(opcode_type, 16#0A#),
      1477 => to_slv(opcode_type, 16#0B#),
      1478 => to_slv(opcode_type, 16#02#),
      1479 => to_slv(opcode_type, 16#0E#),
      1480 => to_slv(opcode_type, 16#11#),
      1481 => to_slv(opcode_type, 16#0C#),
      1482 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#05#),
      1505 => to_slv(opcode_type, 16#07#),
      1506 => to_slv(opcode_type, 16#02#),
      1507 => to_slv(opcode_type, 16#03#),
      1508 => to_slv(opcode_type, 16#78#),
      1509 => to_slv(opcode_type, 16#06#),
      1510 => to_slv(opcode_type, 16#09#),
      1511 => to_slv(opcode_type, 16#59#),
      1512 => to_slv(opcode_type, 16#0F#),
      1513 => to_slv(opcode_type, 16#10#),
      1514 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#06#),
      1537 => to_slv(opcode_type, 16#06#),
      1538 => to_slv(opcode_type, 16#09#),
      1539 => to_slv(opcode_type, 16#07#),
      1540 => to_slv(opcode_type, 16#EB#),
      1541 => to_slv(opcode_type, 16#10#),
      1542 => to_slv(opcode_type, 16#02#),
      1543 => to_slv(opcode_type, 16#11#),
      1544 => to_slv(opcode_type, 16#0F#),
      1545 => to_slv(opcode_type, 16#0C#),
      1546 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#01#),
      1569 => to_slv(opcode_type, 16#08#),
      1570 => to_slv(opcode_type, 16#08#),
      1571 => to_slv(opcode_type, 16#02#),
      1572 => to_slv(opcode_type, 16#0B#),
      1573 => to_slv(opcode_type, 16#08#),
      1574 => to_slv(opcode_type, 16#D7#),
      1575 => to_slv(opcode_type, 16#0E#),
      1576 => to_slv(opcode_type, 16#05#),
      1577 => to_slv(opcode_type, 16#0B#),
      1578 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#05#),
      1601 => to_slv(opcode_type, 16#07#),
      1602 => to_slv(opcode_type, 16#01#),
      1603 => to_slv(opcode_type, 16#09#),
      1604 => to_slv(opcode_type, 16#0C#),
      1605 => to_slv(opcode_type, 16#10#),
      1606 => to_slv(opcode_type, 16#08#),
      1607 => to_slv(opcode_type, 16#04#),
      1608 => to_slv(opcode_type, 16#0E#),
      1609 => to_slv(opcode_type, 16#0E#),
      1610 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#08#),
      1633 => to_slv(opcode_type, 16#07#),
      1634 => to_slv(opcode_type, 16#01#),
      1635 => to_slv(opcode_type, 16#03#),
      1636 => to_slv(opcode_type, 16#11#),
      1637 => to_slv(opcode_type, 16#07#),
      1638 => to_slv(opcode_type, 16#01#),
      1639 => to_slv(opcode_type, 16#0F#),
      1640 => to_slv(opcode_type, 16#0B#),
      1641 => to_slv(opcode_type, 16#0C#),
      1642 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#04#),
      1665 => to_slv(opcode_type, 16#08#),
      1666 => to_slv(opcode_type, 16#06#),
      1667 => to_slv(opcode_type, 16#02#),
      1668 => to_slv(opcode_type, 16#0C#),
      1669 => to_slv(opcode_type, 16#04#),
      1670 => to_slv(opcode_type, 16#0C#),
      1671 => to_slv(opcode_type, 16#09#),
      1672 => to_slv(opcode_type, 16#0F#),
      1673 => to_slv(opcode_type, 16#0B#),
      1674 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#04#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#01#),
      1699 => to_slv(opcode_type, 16#08#),
      1700 => to_slv(opcode_type, 16#0E#),
      1701 => to_slv(opcode_type, 16#0A#),
      1702 => to_slv(opcode_type, 16#05#),
      1703 => to_slv(opcode_type, 16#07#),
      1704 => to_slv(opcode_type, 16#0B#),
      1705 => to_slv(opcode_type, 16#0E#),
      1706 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#04#),
      1729 => to_slv(opcode_type, 16#08#),
      1730 => to_slv(opcode_type, 16#01#),
      1731 => to_slv(opcode_type, 16#03#),
      1732 => to_slv(opcode_type, 16#0C#),
      1733 => to_slv(opcode_type, 16#07#),
      1734 => to_slv(opcode_type, 16#06#),
      1735 => to_slv(opcode_type, 16#0F#),
      1736 => to_slv(opcode_type, 16#0D#),
      1737 => to_slv(opcode_type, 16#11#),
      1738 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#08#),
      1761 => to_slv(opcode_type, 16#07#),
      1762 => to_slv(opcode_type, 16#05#),
      1763 => to_slv(opcode_type, 16#04#),
      1764 => to_slv(opcode_type, 16#10#),
      1765 => to_slv(opcode_type, 16#01#),
      1766 => to_slv(opcode_type, 16#01#),
      1767 => to_slv(opcode_type, 16#11#),
      1768 => to_slv(opcode_type, 16#03#),
      1769 => to_slv(opcode_type, 16#0E#),
      1770 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#01#),
      1793 => to_slv(opcode_type, 16#07#),
      1794 => to_slv(opcode_type, 16#04#),
      1795 => to_slv(opcode_type, 16#01#),
      1796 => to_slv(opcode_type, 16#0F#),
      1797 => to_slv(opcode_type, 16#07#),
      1798 => to_slv(opcode_type, 16#03#),
      1799 => to_slv(opcode_type, 16#0C#),
      1800 => to_slv(opcode_type, 16#03#),
      1801 => to_slv(opcode_type, 16#10#),
      1802 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#09#),
      1825 => to_slv(opcode_type, 16#04#),
      1826 => to_slv(opcode_type, 16#03#),
      1827 => to_slv(opcode_type, 16#02#),
      1828 => to_slv(opcode_type, 16#E3#),
      1829 => to_slv(opcode_type, 16#07#),
      1830 => to_slv(opcode_type, 16#06#),
      1831 => to_slv(opcode_type, 16#0C#),
      1832 => to_slv(opcode_type, 16#0C#),
      1833 => to_slv(opcode_type, 16#0D#),
      1834 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#01#),
      1857 => to_slv(opcode_type, 16#07#),
      1858 => to_slv(opcode_type, 16#02#),
      1859 => to_slv(opcode_type, 16#08#),
      1860 => to_slv(opcode_type, 16#0F#),
      1861 => to_slv(opcode_type, 16#0D#),
      1862 => to_slv(opcode_type, 16#02#),
      1863 => to_slv(opcode_type, 16#07#),
      1864 => to_slv(opcode_type, 16#0A#),
      1865 => to_slv(opcode_type, 16#0C#),
      1866 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#02#),
      1889 => to_slv(opcode_type, 16#06#),
      1890 => to_slv(opcode_type, 16#07#),
      1891 => to_slv(opcode_type, 16#07#),
      1892 => to_slv(opcode_type, 16#DE#),
      1893 => to_slv(opcode_type, 16#0B#),
      1894 => to_slv(opcode_type, 16#05#),
      1895 => to_slv(opcode_type, 16#0A#),
      1896 => to_slv(opcode_type, 16#04#),
      1897 => to_slv(opcode_type, 16#0D#),
      1898 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#03#),
      1921 => to_slv(opcode_type, 16#07#),
      1922 => to_slv(opcode_type, 16#02#),
      1923 => to_slv(opcode_type, 16#05#),
      1924 => to_slv(opcode_type, 16#0F#),
      1925 => to_slv(opcode_type, 16#08#),
      1926 => to_slv(opcode_type, 16#09#),
      1927 => to_slv(opcode_type, 16#0B#),
      1928 => to_slv(opcode_type, 16#EE#),
      1929 => to_slv(opcode_type, 16#0E#),
      1930 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#03#),
      1953 => to_slv(opcode_type, 16#08#),
      1954 => to_slv(opcode_type, 16#04#),
      1955 => to_slv(opcode_type, 16#04#),
      1956 => to_slv(opcode_type, 16#0D#),
      1957 => to_slv(opcode_type, 16#09#),
      1958 => to_slv(opcode_type, 16#05#),
      1959 => to_slv(opcode_type, 16#D7#),
      1960 => to_slv(opcode_type, 16#03#),
      1961 => to_slv(opcode_type, 16#0E#),
      1962 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#03#),
      1985 => to_slv(opcode_type, 16#09#),
      1986 => to_slv(opcode_type, 16#08#),
      1987 => to_slv(opcode_type, 16#07#),
      1988 => to_slv(opcode_type, 16#C0#),
      1989 => to_slv(opcode_type, 16#10#),
      1990 => to_slv(opcode_type, 16#03#),
      1991 => to_slv(opcode_type, 16#0E#),
      1992 => to_slv(opcode_type, 16#01#),
      1993 => to_slv(opcode_type, 16#0D#),
      1994 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#01#),
      2017 => to_slv(opcode_type, 16#07#),
      2018 => to_slv(opcode_type, 16#04#),
      2019 => to_slv(opcode_type, 16#06#),
      2020 => to_slv(opcode_type, 16#0B#),
      2021 => to_slv(opcode_type, 16#11#),
      2022 => to_slv(opcode_type, 16#09#),
      2023 => to_slv(opcode_type, 16#02#),
      2024 => to_slv(opcode_type, 16#0C#),
      2025 => to_slv(opcode_type, 16#0D#),
      2026 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#03#),
      2049 => to_slv(opcode_type, 16#09#),
      2050 => to_slv(opcode_type, 16#08#),
      2051 => to_slv(opcode_type, 16#01#),
      2052 => to_slv(opcode_type, 16#0F#),
      2053 => to_slv(opcode_type, 16#02#),
      2054 => to_slv(opcode_type, 16#0D#),
      2055 => to_slv(opcode_type, 16#02#),
      2056 => to_slv(opcode_type, 16#01#),
      2057 => to_slv(opcode_type, 16#0E#),
      2058 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#08#),
      2081 => to_slv(opcode_type, 16#03#),
      2082 => to_slv(opcode_type, 16#04#),
      2083 => to_slv(opcode_type, 16#07#),
      2084 => to_slv(opcode_type, 16#10#),
      2085 => to_slv(opcode_type, 16#0C#),
      2086 => to_slv(opcode_type, 16#03#),
      2087 => to_slv(opcode_type, 16#08#),
      2088 => to_slv(opcode_type, 16#0C#),
      2089 => to_slv(opcode_type, 16#0A#),
      2090 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#09#),
      2113 => to_slv(opcode_type, 16#05#),
      2114 => to_slv(opcode_type, 16#08#),
      2115 => to_slv(opcode_type, 16#07#),
      2116 => to_slv(opcode_type, 16#0C#),
      2117 => to_slv(opcode_type, 16#10#),
      2118 => to_slv(opcode_type, 16#09#),
      2119 => to_slv(opcode_type, 16#10#),
      2120 => to_slv(opcode_type, 16#11#),
      2121 => to_slv(opcode_type, 16#0F#),
      2122 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#08#),
      2145 => to_slv(opcode_type, 16#06#),
      2146 => to_slv(opcode_type, 16#07#),
      2147 => to_slv(opcode_type, 16#04#),
      2148 => to_slv(opcode_type, 16#10#),
      2149 => to_slv(opcode_type, 16#03#),
      2150 => to_slv(opcode_type, 16#0C#),
      2151 => to_slv(opcode_type, 16#01#),
      2152 => to_slv(opcode_type, 16#0B#),
      2153 => to_slv(opcode_type, 16#0A#),
      2154 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#07#),
      2177 => to_slv(opcode_type, 16#02#),
      2178 => to_slv(opcode_type, 16#03#),
      2179 => to_slv(opcode_type, 16#01#),
      2180 => to_slv(opcode_type, 16#0A#),
      2181 => to_slv(opcode_type, 16#07#),
      2182 => to_slv(opcode_type, 16#04#),
      2183 => to_slv(opcode_type, 16#02#),
      2184 => to_slv(opcode_type, 16#0A#),
      2185 => to_slv(opcode_type, 16#11#),
      2186 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#05#),
      2209 => to_slv(opcode_type, 16#08#),
      2210 => to_slv(opcode_type, 16#09#),
      2211 => to_slv(opcode_type, 16#02#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#02#),
      2214 => to_slv(opcode_type, 16#10#),
      2215 => to_slv(opcode_type, 16#06#),
      2216 => to_slv(opcode_type, 16#0D#),
      2217 => to_slv(opcode_type, 16#0B#),
      2218 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#05#),
      2241 => to_slv(opcode_type, 16#06#),
      2242 => to_slv(opcode_type, 16#09#),
      2243 => to_slv(opcode_type, 16#06#),
      2244 => to_slv(opcode_type, 16#0E#),
      2245 => to_slv(opcode_type, 16#10#),
      2246 => to_slv(opcode_type, 16#08#),
      2247 => to_slv(opcode_type, 16#0B#),
      2248 => to_slv(opcode_type, 16#0A#),
      2249 => to_slv(opcode_type, 16#0D#),
      2250 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#08#),
      2273 => to_slv(opcode_type, 16#05#),
      2274 => to_slv(opcode_type, 16#09#),
      2275 => to_slv(opcode_type, 16#09#),
      2276 => to_slv(opcode_type, 16#0F#),
      2277 => to_slv(opcode_type, 16#0F#),
      2278 => to_slv(opcode_type, 16#06#),
      2279 => to_slv(opcode_type, 16#0A#),
      2280 => to_slv(opcode_type, 16#0C#),
      2281 => to_slv(opcode_type, 16#A3#),
      2282 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#07#),
      2305 => to_slv(opcode_type, 16#05#),
      2306 => to_slv(opcode_type, 16#04#),
      2307 => to_slv(opcode_type, 16#07#),
      2308 => to_slv(opcode_type, 16#10#),
      2309 => to_slv(opcode_type, 16#FB#),
      2310 => to_slv(opcode_type, 16#07#),
      2311 => to_slv(opcode_type, 16#05#),
      2312 => to_slv(opcode_type, 16#0C#),
      2313 => to_slv(opcode_type, 16#10#),
      2314 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#01#),
      2337 => to_slv(opcode_type, 16#09#),
      2338 => to_slv(opcode_type, 16#09#),
      2339 => to_slv(opcode_type, 16#02#),
      2340 => to_slv(opcode_type, 16#0E#),
      2341 => to_slv(opcode_type, 16#08#),
      2342 => to_slv(opcode_type, 16#F4#),
      2343 => to_slv(opcode_type, 16#0E#),
      2344 => to_slv(opcode_type, 16#03#),
      2345 => to_slv(opcode_type, 16#0B#),
      2346 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#01#),
      2369 => to_slv(opcode_type, 16#06#),
      2370 => to_slv(opcode_type, 16#03#),
      2371 => to_slv(opcode_type, 16#04#),
      2372 => to_slv(opcode_type, 16#0F#),
      2373 => to_slv(opcode_type, 16#06#),
      2374 => to_slv(opcode_type, 16#05#),
      2375 => to_slv(opcode_type, 16#0F#),
      2376 => to_slv(opcode_type, 16#05#),
      2377 => to_slv(opcode_type, 16#0D#),
      2378 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#02#),
      2402 => to_slv(opcode_type, 16#06#),
      2403 => to_slv(opcode_type, 16#09#),
      2404 => to_slv(opcode_type, 16#0C#),
      2405 => to_slv(opcode_type, 16#0B#),
      2406 => to_slv(opcode_type, 16#02#),
      2407 => to_slv(opcode_type, 16#0B#),
      2408 => to_slv(opcode_type, 16#04#),
      2409 => to_slv(opcode_type, 16#3F#),
      2410 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#05#),
      2433 => to_slv(opcode_type, 16#07#),
      2434 => to_slv(opcode_type, 16#02#),
      2435 => to_slv(opcode_type, 16#03#),
      2436 => to_slv(opcode_type, 16#0B#),
      2437 => to_slv(opcode_type, 16#06#),
      2438 => to_slv(opcode_type, 16#02#),
      2439 => to_slv(opcode_type, 16#10#),
      2440 => to_slv(opcode_type, 16#02#),
      2441 => to_slv(opcode_type, 16#0F#),
      2442 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#09#),
      2465 => to_slv(opcode_type, 16#01#),
      2466 => to_slv(opcode_type, 16#08#),
      2467 => to_slv(opcode_type, 16#02#),
      2468 => to_slv(opcode_type, 16#10#),
      2469 => to_slv(opcode_type, 16#07#),
      2470 => to_slv(opcode_type, 16#2F#),
      2471 => to_slv(opcode_type, 16#10#),
      2472 => to_slv(opcode_type, 16#04#),
      2473 => to_slv(opcode_type, 16#0F#),
      2474 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#01#),
      2497 => to_slv(opcode_type, 16#06#),
      2498 => to_slv(opcode_type, 16#07#),
      2499 => to_slv(opcode_type, 16#09#),
      2500 => to_slv(opcode_type, 16#0B#),
      2501 => to_slv(opcode_type, 16#0E#),
      2502 => to_slv(opcode_type, 16#06#),
      2503 => to_slv(opcode_type, 16#0B#),
      2504 => to_slv(opcode_type, 16#0F#),
      2505 => to_slv(opcode_type, 16#10#),
      2506 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#01#),
      2529 => to_slv(opcode_type, 16#08#),
      2530 => to_slv(opcode_type, 16#09#),
      2531 => to_slv(opcode_type, 16#04#),
      2532 => to_slv(opcode_type, 16#0C#),
      2533 => to_slv(opcode_type, 16#05#),
      2534 => to_slv(opcode_type, 16#11#),
      2535 => to_slv(opcode_type, 16#03#),
      2536 => to_slv(opcode_type, 16#03#),
      2537 => to_slv(opcode_type, 16#10#),
      2538 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#03#),
      2561 => to_slv(opcode_type, 16#07#),
      2562 => to_slv(opcode_type, 16#05#),
      2563 => to_slv(opcode_type, 16#03#),
      2564 => to_slv(opcode_type, 16#10#),
      2565 => to_slv(opcode_type, 16#08#),
      2566 => to_slv(opcode_type, 16#06#),
      2567 => to_slv(opcode_type, 16#0F#),
      2568 => to_slv(opcode_type, 16#11#),
      2569 => to_slv(opcode_type, 16#0B#),
      2570 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#04#),
      2593 => to_slv(opcode_type, 16#06#),
      2594 => to_slv(opcode_type, 16#04#),
      2595 => to_slv(opcode_type, 16#06#),
      2596 => to_slv(opcode_type, 16#11#),
      2597 => to_slv(opcode_type, 16#0F#),
      2598 => to_slv(opcode_type, 16#03#),
      2599 => to_slv(opcode_type, 16#08#),
      2600 => to_slv(opcode_type, 16#0C#),
      2601 => to_slv(opcode_type, 16#0B#),
      2602 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#06#),
      2625 => to_slv(opcode_type, 16#08#),
      2626 => to_slv(opcode_type, 16#06#),
      2627 => to_slv(opcode_type, 16#08#),
      2628 => to_slv(opcode_type, 16#0C#),
      2629 => to_slv(opcode_type, 16#0B#),
      2630 => to_slv(opcode_type, 16#04#),
      2631 => to_slv(opcode_type, 16#0C#),
      2632 => to_slv(opcode_type, 16#0A#),
      2633 => to_slv(opcode_type, 16#0D#),
      2634 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#06#),
      2657 => to_slv(opcode_type, 16#04#),
      2658 => to_slv(opcode_type, 16#08#),
      2659 => to_slv(opcode_type, 16#03#),
      2660 => to_slv(opcode_type, 16#0A#),
      2661 => to_slv(opcode_type, 16#08#),
      2662 => to_slv(opcode_type, 16#11#),
      2663 => to_slv(opcode_type, 16#0C#),
      2664 => to_slv(opcode_type, 16#05#),
      2665 => to_slv(opcode_type, 16#10#),
      2666 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#09#),
      2689 => to_slv(opcode_type, 16#05#),
      2690 => to_slv(opcode_type, 16#06#),
      2691 => to_slv(opcode_type, 16#06#),
      2692 => to_slv(opcode_type, 16#11#),
      2693 => to_slv(opcode_type, 16#10#),
      2694 => to_slv(opcode_type, 16#01#),
      2695 => to_slv(opcode_type, 16#0C#),
      2696 => to_slv(opcode_type, 16#01#),
      2697 => to_slv(opcode_type, 16#10#),
      2698 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#07#),
      2721 => to_slv(opcode_type, 16#05#),
      2722 => to_slv(opcode_type, 16#06#),
      2723 => to_slv(opcode_type, 16#09#),
      2724 => to_slv(opcode_type, 16#2E#),
      2725 => to_slv(opcode_type, 16#0A#),
      2726 => to_slv(opcode_type, 16#06#),
      2727 => to_slv(opcode_type, 16#11#),
      2728 => to_slv(opcode_type, 16#0F#),
      2729 => to_slv(opcode_type, 16#8F#),
      2730 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#09#),
      2753 => to_slv(opcode_type, 16#06#),
      2754 => to_slv(opcode_type, 16#06#),
      2755 => to_slv(opcode_type, 16#08#),
      2756 => to_slv(opcode_type, 16#AC#),
      2757 => to_slv(opcode_type, 16#C5#),
      2758 => to_slv(opcode_type, 16#04#),
      2759 => to_slv(opcode_type, 16#0E#),
      2760 => to_slv(opcode_type, 16#24#),
      2761 => to_slv(opcode_type, 16#11#),
      2762 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#07#),
      2785 => to_slv(opcode_type, 16#05#),
      2786 => to_slv(opcode_type, 16#09#),
      2787 => to_slv(opcode_type, 16#06#),
      2788 => to_slv(opcode_type, 16#0C#),
      2789 => to_slv(opcode_type, 16#0C#),
      2790 => to_slv(opcode_type, 16#05#),
      2791 => to_slv(opcode_type, 16#0E#),
      2792 => to_slv(opcode_type, 16#03#),
      2793 => to_slv(opcode_type, 16#11#),
      2794 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#07#),
      2817 => to_slv(opcode_type, 16#03#),
      2818 => to_slv(opcode_type, 16#07#),
      2819 => to_slv(opcode_type, 16#06#),
      2820 => to_slv(opcode_type, 16#0A#),
      2821 => to_slv(opcode_type, 16#31#),
      2822 => to_slv(opcode_type, 16#09#),
      2823 => to_slv(opcode_type, 16#0E#),
      2824 => to_slv(opcode_type, 16#0B#),
      2825 => to_slv(opcode_type, 16#DA#),
      2826 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#06#),
      2849 => to_slv(opcode_type, 16#06#),
      2850 => to_slv(opcode_type, 16#01#),
      2851 => to_slv(opcode_type, 16#04#),
      2852 => to_slv(opcode_type, 16#0A#),
      2853 => to_slv(opcode_type, 16#02#),
      2854 => to_slv(opcode_type, 16#02#),
      2855 => to_slv(opcode_type, 16#0E#),
      2856 => to_slv(opcode_type, 16#03#),
      2857 => to_slv(opcode_type, 16#10#),
      2858 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#05#),
      2881 => to_slv(opcode_type, 16#09#),
      2882 => to_slv(opcode_type, 16#02#),
      2883 => to_slv(opcode_type, 16#05#),
      2884 => to_slv(opcode_type, 16#10#),
      2885 => to_slv(opcode_type, 16#08#),
      2886 => to_slv(opcode_type, 16#09#),
      2887 => to_slv(opcode_type, 16#10#),
      2888 => to_slv(opcode_type, 16#0C#),
      2889 => to_slv(opcode_type, 16#68#),
      2890 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#03#),
      2913 => to_slv(opcode_type, 16#08#),
      2914 => to_slv(opcode_type, 16#01#),
      2915 => to_slv(opcode_type, 16#03#),
      2916 => to_slv(opcode_type, 16#0F#),
      2917 => to_slv(opcode_type, 16#09#),
      2918 => to_slv(opcode_type, 16#07#),
      2919 => to_slv(opcode_type, 16#10#),
      2920 => to_slv(opcode_type, 16#11#),
      2921 => to_slv(opcode_type, 16#0B#),
      2922 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#01#),
      2945 => to_slv(opcode_type, 16#09#),
      2946 => to_slv(opcode_type, 16#04#),
      2947 => to_slv(opcode_type, 16#03#),
      2948 => to_slv(opcode_type, 16#0F#),
      2949 => to_slv(opcode_type, 16#07#),
      2950 => to_slv(opcode_type, 16#08#),
      2951 => to_slv(opcode_type, 16#0B#),
      2952 => to_slv(opcode_type, 16#0F#),
      2953 => to_slv(opcode_type, 16#0B#),
      2954 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#03#),
      2977 => to_slv(opcode_type, 16#06#),
      2978 => to_slv(opcode_type, 16#06#),
      2979 => to_slv(opcode_type, 16#08#),
      2980 => to_slv(opcode_type, 16#0B#),
      2981 => to_slv(opcode_type, 16#0A#),
      2982 => to_slv(opcode_type, 16#06#),
      2983 => to_slv(opcode_type, 16#10#),
      2984 => to_slv(opcode_type, 16#0F#),
      2985 => to_slv(opcode_type, 16#0D#),
      2986 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#08#),
      3009 => to_slv(opcode_type, 16#03#),
      3010 => to_slv(opcode_type, 16#07#),
      3011 => to_slv(opcode_type, 16#03#),
      3012 => to_slv(opcode_type, 16#0F#),
      3013 => to_slv(opcode_type, 16#03#),
      3014 => to_slv(opcode_type, 16#0B#),
      3015 => to_slv(opcode_type, 16#07#),
      3016 => to_slv(opcode_type, 16#0B#),
      3017 => to_slv(opcode_type, 16#10#),
      3018 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#02#),
      3041 => to_slv(opcode_type, 16#09#),
      3042 => to_slv(opcode_type, 16#07#),
      3043 => to_slv(opcode_type, 16#02#),
      3044 => to_slv(opcode_type, 16#0C#),
      3045 => to_slv(opcode_type, 16#03#),
      3046 => to_slv(opcode_type, 16#0C#),
      3047 => to_slv(opcode_type, 16#02#),
      3048 => to_slv(opcode_type, 16#05#),
      3049 => to_slv(opcode_type, 16#0F#),
      3050 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#09#),
      3073 => to_slv(opcode_type, 16#09#),
      3074 => to_slv(opcode_type, 16#03#),
      3075 => to_slv(opcode_type, 16#05#),
      3076 => to_slv(opcode_type, 16#8E#),
      3077 => to_slv(opcode_type, 16#03#),
      3078 => to_slv(opcode_type, 16#08#),
      3079 => to_slv(opcode_type, 16#0D#),
      3080 => to_slv(opcode_type, 16#10#),
      3081 => to_slv(opcode_type, 16#10#),
      3082 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#05#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#08#),
      3107 => to_slv(opcode_type, 16#09#),
      3108 => to_slv(opcode_type, 16#11#),
      3109 => to_slv(opcode_type, 16#0D#),
      3110 => to_slv(opcode_type, 16#07#),
      3111 => to_slv(opcode_type, 16#0C#),
      3112 => to_slv(opcode_type, 16#0D#),
      3113 => to_slv(opcode_type, 16#0E#),
      3114 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#07#),
      3137 => to_slv(opcode_type, 16#09#),
      3138 => to_slv(opcode_type, 16#08#),
      3139 => to_slv(opcode_type, 16#08#),
      3140 => to_slv(opcode_type, 16#B4#),
      3141 => to_slv(opcode_type, 16#0F#),
      3142 => to_slv(opcode_type, 16#05#),
      3143 => to_slv(opcode_type, 16#0A#),
      3144 => to_slv(opcode_type, 16#0F#),
      3145 => to_slv(opcode_type, 16#0C#),
      3146 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#07#),
      3169 => to_slv(opcode_type, 16#04#),
      3170 => to_slv(opcode_type, 16#02#),
      3171 => to_slv(opcode_type, 16#02#),
      3172 => to_slv(opcode_type, 16#0D#),
      3173 => to_slv(opcode_type, 16#01#),
      3174 => to_slv(opcode_type, 16#04#),
      3175 => to_slv(opcode_type, 16#06#),
      3176 => to_slv(opcode_type, 16#0E#),
      3177 => to_slv(opcode_type, 16#10#),
      3178 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#07#),
      3201 => to_slv(opcode_type, 16#01#),
      3202 => to_slv(opcode_type, 16#09#),
      3203 => to_slv(opcode_type, 16#08#),
      3204 => to_slv(opcode_type, 16#6F#),
      3205 => to_slv(opcode_type, 16#0D#),
      3206 => to_slv(opcode_type, 16#09#),
      3207 => to_slv(opcode_type, 16#11#),
      3208 => to_slv(opcode_type, 16#0D#),
      3209 => to_slv(opcode_type, 16#0E#),
      3210 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#05#),
      3234 => to_slv(opcode_type, 16#09#),
      3235 => to_slv(opcode_type, 16#06#),
      3236 => to_slv(opcode_type, 16#0C#),
      3237 => to_slv(opcode_type, 16#0B#),
      3238 => to_slv(opcode_type, 16#02#),
      3239 => to_slv(opcode_type, 16#10#),
      3240 => to_slv(opcode_type, 16#05#),
      3241 => to_slv(opcode_type, 16#11#),
      3242 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#09#),
      3265 => to_slv(opcode_type, 16#08#),
      3266 => to_slv(opcode_type, 16#01#),
      3267 => to_slv(opcode_type, 16#01#),
      3268 => to_slv(opcode_type, 16#0D#),
      3269 => to_slv(opcode_type, 16#03#),
      3270 => to_slv(opcode_type, 16#05#),
      3271 => to_slv(opcode_type, 16#BC#),
      3272 => to_slv(opcode_type, 16#01#),
      3273 => to_slv(opcode_type, 16#BF#),
      3274 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#08#),
      3297 => to_slv(opcode_type, 16#05#),
      3298 => to_slv(opcode_type, 16#02#),
      3299 => to_slv(opcode_type, 16#05#),
      3300 => to_slv(opcode_type, 16#0E#),
      3301 => to_slv(opcode_type, 16#09#),
      3302 => to_slv(opcode_type, 16#08#),
      3303 => to_slv(opcode_type, 16#0C#),
      3304 => to_slv(opcode_type, 16#10#),
      3305 => to_slv(opcode_type, 16#46#),
      3306 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#04#),
      3329 => to_slv(opcode_type, 16#08#),
      3330 => to_slv(opcode_type, 16#09#),
      3331 => to_slv(opcode_type, 16#05#),
      3332 => to_slv(opcode_type, 16#0E#),
      3333 => to_slv(opcode_type, 16#09#),
      3334 => to_slv(opcode_type, 16#AE#),
      3335 => to_slv(opcode_type, 16#0A#),
      3336 => to_slv(opcode_type, 16#04#),
      3337 => to_slv(opcode_type, 16#10#),
      3338 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#03#),
      3361 => to_slv(opcode_type, 16#06#),
      3362 => to_slv(opcode_type, 16#07#),
      3363 => to_slv(opcode_type, 16#05#),
      3364 => to_slv(opcode_type, 16#0E#),
      3365 => to_slv(opcode_type, 16#09#),
      3366 => to_slv(opcode_type, 16#0C#),
      3367 => to_slv(opcode_type, 16#0E#),
      3368 => to_slv(opcode_type, 16#03#),
      3369 => to_slv(opcode_type, 16#0A#),
      3370 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#09#),
      3393 => to_slv(opcode_type, 16#02#),
      3394 => to_slv(opcode_type, 16#04#),
      3395 => to_slv(opcode_type, 16#09#),
      3396 => to_slv(opcode_type, 16#0B#),
      3397 => to_slv(opcode_type, 16#0B#),
      3398 => to_slv(opcode_type, 16#03#),
      3399 => to_slv(opcode_type, 16#04#),
      3400 => to_slv(opcode_type, 16#01#),
      3401 => to_slv(opcode_type, 16#0B#),
      3402 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#02#),
      3425 => to_slv(opcode_type, 16#08#),
      3426 => to_slv(opcode_type, 16#05#),
      3427 => to_slv(opcode_type, 16#08#),
      3428 => to_slv(opcode_type, 16#0D#),
      3429 => to_slv(opcode_type, 16#69#),
      3430 => to_slv(opcode_type, 16#03#),
      3431 => to_slv(opcode_type, 16#06#),
      3432 => to_slv(opcode_type, 16#0E#),
      3433 => to_slv(opcode_type, 16#11#),
      3434 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#09#),
      3457 => to_slv(opcode_type, 16#08#),
      3458 => to_slv(opcode_type, 16#01#),
      3459 => to_slv(opcode_type, 16#02#),
      3460 => to_slv(opcode_type, 16#0F#),
      3461 => to_slv(opcode_type, 16#09#),
      3462 => to_slv(opcode_type, 16#04#),
      3463 => to_slv(opcode_type, 16#10#),
      3464 => to_slv(opcode_type, 16#0C#),
      3465 => to_slv(opcode_type, 16#0E#),
      3466 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#09#),
      3489 => to_slv(opcode_type, 16#03#),
      3490 => to_slv(opcode_type, 16#06#),
      3491 => to_slv(opcode_type, 16#07#),
      3492 => to_slv(opcode_type, 16#0C#),
      3493 => to_slv(opcode_type, 16#0F#),
      3494 => to_slv(opcode_type, 16#08#),
      3495 => to_slv(opcode_type, 16#10#),
      3496 => to_slv(opcode_type, 16#0E#),
      3497 => to_slv(opcode_type, 16#6B#),
      3498 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#04#),
      3521 => to_slv(opcode_type, 16#07#),
      3522 => to_slv(opcode_type, 16#02#),
      3523 => to_slv(opcode_type, 16#07#),
      3524 => to_slv(opcode_type, 16#0F#),
      3525 => to_slv(opcode_type, 16#0A#),
      3526 => to_slv(opcode_type, 16#04#),
      3527 => to_slv(opcode_type, 16#08#),
      3528 => to_slv(opcode_type, 16#10#),
      3529 => to_slv(opcode_type, 16#11#),
      3530 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#02#),
      3553 => to_slv(opcode_type, 16#06#),
      3554 => to_slv(opcode_type, 16#05#),
      3555 => to_slv(opcode_type, 16#02#),
      3556 => to_slv(opcode_type, 16#0E#),
      3557 => to_slv(opcode_type, 16#09#),
      3558 => to_slv(opcode_type, 16#04#),
      3559 => to_slv(opcode_type, 16#0C#),
      3560 => to_slv(opcode_type, 16#02#),
      3561 => to_slv(opcode_type, 16#F9#),
      3562 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#09#),
      3585 => to_slv(opcode_type, 16#05#),
      3586 => to_slv(opcode_type, 16#04#),
      3587 => to_slv(opcode_type, 16#03#),
      3588 => to_slv(opcode_type, 16#0B#),
      3589 => to_slv(opcode_type, 16#05#),
      3590 => to_slv(opcode_type, 16#08#),
      3591 => to_slv(opcode_type, 16#05#),
      3592 => to_slv(opcode_type, 16#0C#),
      3593 => to_slv(opcode_type, 16#0F#),
      3594 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#06#),
      3617 => to_slv(opcode_type, 16#02#),
      3618 => to_slv(opcode_type, 16#05#),
      3619 => to_slv(opcode_type, 16#08#),
      3620 => to_slv(opcode_type, 16#0D#),
      3621 => to_slv(opcode_type, 16#98#),
      3622 => to_slv(opcode_type, 16#06#),
      3623 => to_slv(opcode_type, 16#02#),
      3624 => to_slv(opcode_type, 16#0E#),
      3625 => to_slv(opcode_type, 16#0D#),
      3626 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#06#),
      3649 => to_slv(opcode_type, 16#02#),
      3650 => to_slv(opcode_type, 16#09#),
      3651 => to_slv(opcode_type, 16#01#),
      3652 => to_slv(opcode_type, 16#10#),
      3653 => to_slv(opcode_type, 16#03#),
      3654 => to_slv(opcode_type, 16#0E#),
      3655 => to_slv(opcode_type, 16#06#),
      3656 => to_slv(opcode_type, 16#0A#),
      3657 => to_slv(opcode_type, 16#0B#),
      3658 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#04#),
      3681 => to_slv(opcode_type, 16#07#),
      3682 => to_slv(opcode_type, 16#09#),
      3683 => to_slv(opcode_type, 16#09#),
      3684 => to_slv(opcode_type, 16#11#),
      3685 => to_slv(opcode_type, 16#11#),
      3686 => to_slv(opcode_type, 16#02#),
      3687 => to_slv(opcode_type, 16#0D#),
      3688 => to_slv(opcode_type, 16#03#),
      3689 => to_slv(opcode_type, 16#0A#),
      3690 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#01#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#03#),
      3715 => to_slv(opcode_type, 16#07#),
      3716 => to_slv(opcode_type, 16#0D#),
      3717 => to_slv(opcode_type, 16#0E#),
      3718 => to_slv(opcode_type, 16#07#),
      3719 => to_slv(opcode_type, 16#02#),
      3720 => to_slv(opcode_type, 16#0C#),
      3721 => to_slv(opcode_type, 16#0A#),
      3722 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#09#),
      3745 => to_slv(opcode_type, 16#07#),
      3746 => to_slv(opcode_type, 16#03#),
      3747 => to_slv(opcode_type, 16#01#),
      3748 => to_slv(opcode_type, 16#0C#),
      3749 => to_slv(opcode_type, 16#02#),
      3750 => to_slv(opcode_type, 16#04#),
      3751 => to_slv(opcode_type, 16#11#),
      3752 => to_slv(opcode_type, 16#02#),
      3753 => to_slv(opcode_type, 16#10#),
      3754 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#04#),
      3777 => to_slv(opcode_type, 16#08#),
      3778 => to_slv(opcode_type, 16#01#),
      3779 => to_slv(opcode_type, 16#04#),
      3780 => to_slv(opcode_type, 16#0E#),
      3781 => to_slv(opcode_type, 16#06#),
      3782 => to_slv(opcode_type, 16#01#),
      3783 => to_slv(opcode_type, 16#EE#),
      3784 => to_slv(opcode_type, 16#04#),
      3785 => to_slv(opcode_type, 16#11#),
      3786 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#03#),
      3809 => to_slv(opcode_type, 16#07#),
      3810 => to_slv(opcode_type, 16#07#),
      3811 => to_slv(opcode_type, 16#05#),
      3812 => to_slv(opcode_type, 16#10#),
      3813 => to_slv(opcode_type, 16#06#),
      3814 => to_slv(opcode_type, 16#0C#),
      3815 => to_slv(opcode_type, 16#0C#),
      3816 => to_slv(opcode_type, 16#03#),
      3817 => to_slv(opcode_type, 16#0E#),
      3818 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#04#),
      3841 => to_slv(opcode_type, 16#07#),
      3842 => to_slv(opcode_type, 16#05#),
      3843 => to_slv(opcode_type, 16#05#),
      3844 => to_slv(opcode_type, 16#0A#),
      3845 => to_slv(opcode_type, 16#08#),
      3846 => to_slv(opcode_type, 16#01#),
      3847 => to_slv(opcode_type, 16#0D#),
      3848 => to_slv(opcode_type, 16#03#),
      3849 => to_slv(opcode_type, 16#0D#),
      3850 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#02#),
      3873 => to_slv(opcode_type, 16#07#),
      3874 => to_slv(opcode_type, 16#06#),
      3875 => to_slv(opcode_type, 16#07#),
      3876 => to_slv(opcode_type, 16#11#),
      3877 => to_slv(opcode_type, 16#0E#),
      3878 => to_slv(opcode_type, 16#03#),
      3879 => to_slv(opcode_type, 16#0D#),
      3880 => to_slv(opcode_type, 16#01#),
      3881 => to_slv(opcode_type, 16#10#),
      3882 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#08#),
      3905 => to_slv(opcode_type, 16#07#),
      3906 => to_slv(opcode_type, 16#05#),
      3907 => to_slv(opcode_type, 16#06#),
      3908 => to_slv(opcode_type, 16#0F#),
      3909 => to_slv(opcode_type, 16#0E#),
      3910 => to_slv(opcode_type, 16#07#),
      3911 => to_slv(opcode_type, 16#0D#),
      3912 => to_slv(opcode_type, 16#10#),
      3913 => to_slv(opcode_type, 16#10#),
      3914 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#01#),
      3937 => to_slv(opcode_type, 16#07#),
      3938 => to_slv(opcode_type, 16#05#),
      3939 => to_slv(opcode_type, 16#08#),
      3940 => to_slv(opcode_type, 16#0D#),
      3941 => to_slv(opcode_type, 16#0E#),
      3942 => to_slv(opcode_type, 16#05#),
      3943 => to_slv(opcode_type, 16#07#),
      3944 => to_slv(opcode_type, 16#10#),
      3945 => to_slv(opcode_type, 16#7D#),
      3946 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#01#),
      3969 => to_slv(opcode_type, 16#09#),
      3970 => to_slv(opcode_type, 16#04#),
      3971 => to_slv(opcode_type, 16#05#),
      3972 => to_slv(opcode_type, 16#11#),
      3973 => to_slv(opcode_type, 16#06#),
      3974 => to_slv(opcode_type, 16#05#),
      3975 => to_slv(opcode_type, 16#0C#),
      3976 => to_slv(opcode_type, 16#04#),
      3977 => to_slv(opcode_type, 16#0A#),
      3978 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#01#),
      4001 => to_slv(opcode_type, 16#09#),
      4002 => to_slv(opcode_type, 16#08#),
      4003 => to_slv(opcode_type, 16#06#),
      4004 => to_slv(opcode_type, 16#5D#),
      4005 => to_slv(opcode_type, 16#E4#),
      4006 => to_slv(opcode_type, 16#09#),
      4007 => to_slv(opcode_type, 16#95#),
      4008 => to_slv(opcode_type, 16#11#),
      4009 => to_slv(opcode_type, 16#99#),
      4010 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#06#),
      4033 => to_slv(opcode_type, 16#07#),
      4034 => to_slv(opcode_type, 16#02#),
      4035 => to_slv(opcode_type, 16#03#),
      4036 => to_slv(opcode_type, 16#11#),
      4037 => to_slv(opcode_type, 16#03#),
      4038 => to_slv(opcode_type, 16#01#),
      4039 => to_slv(opcode_type, 16#69#),
      4040 => to_slv(opcode_type, 16#05#),
      4041 => to_slv(opcode_type, 16#0E#),
      4042 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#08#),
      4065 => to_slv(opcode_type, 16#06#),
      4066 => to_slv(opcode_type, 16#05#),
      4067 => to_slv(opcode_type, 16#09#),
      4068 => to_slv(opcode_type, 16#11#),
      4069 => to_slv(opcode_type, 16#0C#),
      4070 => to_slv(opcode_type, 16#08#),
      4071 => to_slv(opcode_type, 16#11#),
      4072 => to_slv(opcode_type, 16#0F#),
      4073 => to_slv(opcode_type, 16#0D#),
      4074 to 4095 => (others => '0')
  ),

    -- Bin `11`...
    10 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#07#),
      1 => to_slv(opcode_type, 16#02#),
      2 => to_slv(opcode_type, 16#04#),
      3 => to_slv(opcode_type, 16#09#),
      4 => to_slv(opcode_type, 16#0F#),
      5 => to_slv(opcode_type, 16#11#),
      6 => to_slv(opcode_type, 16#09#),
      7 => to_slv(opcode_type, 16#09#),
      8 => to_slv(opcode_type, 16#0D#),
      9 => to_slv(opcode_type, 16#7F#),
      10 => to_slv(opcode_type, 16#0B#),
      11 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#06#),
      33 => to_slv(opcode_type, 16#06#),
      34 => to_slv(opcode_type, 16#06#),
      35 => to_slv(opcode_type, 16#04#),
      36 => to_slv(opcode_type, 16#11#),
      37 => to_slv(opcode_type, 16#08#),
      38 => to_slv(opcode_type, 16#0C#),
      39 => to_slv(opcode_type, 16#11#),
      40 => to_slv(opcode_type, 16#01#),
      41 => to_slv(opcode_type, 16#0C#),
      42 => to_slv(opcode_type, 16#0D#),
      43 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#02#),
      65 => to_slv(opcode_type, 16#08#),
      66 => to_slv(opcode_type, 16#05#),
      67 => to_slv(opcode_type, 16#01#),
      68 => to_slv(opcode_type, 16#0D#),
      69 => to_slv(opcode_type, 16#07#),
      70 => to_slv(opcode_type, 16#09#),
      71 => to_slv(opcode_type, 16#3F#),
      72 => to_slv(opcode_type, 16#11#),
      73 => to_slv(opcode_type, 16#05#),
      74 => to_slv(opcode_type, 16#0C#),
      75 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#08#),
      97 => to_slv(opcode_type, 16#01#),
      98 => to_slv(opcode_type, 16#03#),
      99 => to_slv(opcode_type, 16#04#),
      100 => to_slv(opcode_type, 16#66#),
      101 => to_slv(opcode_type, 16#08#),
      102 => to_slv(opcode_type, 16#06#),
      103 => to_slv(opcode_type, 16#03#),
      104 => to_slv(opcode_type, 16#0D#),
      105 => to_slv(opcode_type, 16#0F#),
      106 => to_slv(opcode_type, 16#0B#),
      107 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#09#),
      129 => to_slv(opcode_type, 16#05#),
      130 => to_slv(opcode_type, 16#09#),
      131 => to_slv(opcode_type, 16#08#),
      132 => to_slv(opcode_type, 16#11#),
      133 => to_slv(opcode_type, 16#0A#),
      134 => to_slv(opcode_type, 16#01#),
      135 => to_slv(opcode_type, 16#56#),
      136 => to_slv(opcode_type, 16#01#),
      137 => to_slv(opcode_type, 16#03#),
      138 => to_slv(opcode_type, 16#0C#),
      139 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#01#),
      161 => to_slv(opcode_type, 16#09#),
      162 => to_slv(opcode_type, 16#08#),
      163 => to_slv(opcode_type, 16#02#),
      164 => to_slv(opcode_type, 16#10#),
      165 => to_slv(opcode_type, 16#01#),
      166 => to_slv(opcode_type, 16#E5#),
      167 => to_slv(opcode_type, 16#01#),
      168 => to_slv(opcode_type, 16#06#),
      169 => to_slv(opcode_type, 16#2B#),
      170 => to_slv(opcode_type, 16#10#),
      171 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#07#),
      193 => to_slv(opcode_type, 16#09#),
      194 => to_slv(opcode_type, 16#01#),
      195 => to_slv(opcode_type, 16#04#),
      196 => to_slv(opcode_type, 16#0C#),
      197 => to_slv(opcode_type, 16#09#),
      198 => to_slv(opcode_type, 16#07#),
      199 => to_slv(opcode_type, 16#0F#),
      200 => to_slv(opcode_type, 16#19#),
      201 => to_slv(opcode_type, 16#0C#),
      202 => to_slv(opcode_type, 16#0F#),
      203 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#03#),
      225 => to_slv(opcode_type, 16#08#),
      226 => to_slv(opcode_type, 16#07#),
      227 => to_slv(opcode_type, 16#09#),
      228 => to_slv(opcode_type, 16#0D#),
      229 => to_slv(opcode_type, 16#0D#),
      230 => to_slv(opcode_type, 16#09#),
      231 => to_slv(opcode_type, 16#0D#),
      232 => to_slv(opcode_type, 16#D8#),
      233 => to_slv(opcode_type, 16#02#),
      234 => to_slv(opcode_type, 16#10#),
      235 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#02#),
      257 => to_slv(opcode_type, 16#09#),
      258 => to_slv(opcode_type, 16#05#),
      259 => to_slv(opcode_type, 16#07#),
      260 => to_slv(opcode_type, 16#0F#),
      261 => to_slv(opcode_type, 16#0B#),
      262 => to_slv(opcode_type, 16#09#),
      263 => to_slv(opcode_type, 16#04#),
      264 => to_slv(opcode_type, 16#11#),
      265 => to_slv(opcode_type, 16#02#),
      266 => to_slv(opcode_type, 16#11#),
      267 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#03#),
      289 => to_slv(opcode_type, 16#08#),
      290 => to_slv(opcode_type, 16#08#),
      291 => to_slv(opcode_type, 16#01#),
      292 => to_slv(opcode_type, 16#10#),
      293 => to_slv(opcode_type, 16#03#),
      294 => to_slv(opcode_type, 16#0F#),
      295 => to_slv(opcode_type, 16#02#),
      296 => to_slv(opcode_type, 16#09#),
      297 => to_slv(opcode_type, 16#0C#),
      298 => to_slv(opcode_type, 16#10#),
      299 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#01#),
      321 => to_slv(opcode_type, 16#07#),
      322 => to_slv(opcode_type, 16#03#),
      323 => to_slv(opcode_type, 16#04#),
      324 => to_slv(opcode_type, 16#0D#),
      325 => to_slv(opcode_type, 16#06#),
      326 => to_slv(opcode_type, 16#06#),
      327 => to_slv(opcode_type, 16#0D#),
      328 => to_slv(opcode_type, 16#11#),
      329 => to_slv(opcode_type, 16#03#),
      330 => to_slv(opcode_type, 16#0C#),
      331 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#07#),
      353 => to_slv(opcode_type, 16#08#),
      354 => to_slv(opcode_type, 16#02#),
      355 => to_slv(opcode_type, 16#08#),
      356 => to_slv(opcode_type, 16#0C#),
      357 => to_slv(opcode_type, 16#0A#),
      358 => to_slv(opcode_type, 16#08#),
      359 => to_slv(opcode_type, 16#05#),
      360 => to_slv(opcode_type, 16#0D#),
      361 => to_slv(opcode_type, 16#E1#),
      362 => to_slv(opcode_type, 16#0B#),
      363 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#02#),
      385 => to_slv(opcode_type, 16#07#),
      386 => to_slv(opcode_type, 16#05#),
      387 => to_slv(opcode_type, 16#05#),
      388 => to_slv(opcode_type, 16#10#),
      389 => to_slv(opcode_type, 16#07#),
      390 => to_slv(opcode_type, 16#05#),
      391 => to_slv(opcode_type, 16#0C#),
      392 => to_slv(opcode_type, 16#09#),
      393 => to_slv(opcode_type, 16#0D#),
      394 => to_slv(opcode_type, 16#10#),
      395 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#03#),
      417 => to_slv(opcode_type, 16#06#),
      418 => to_slv(opcode_type, 16#07#),
      419 => to_slv(opcode_type, 16#06#),
      420 => to_slv(opcode_type, 16#10#),
      421 => to_slv(opcode_type, 16#0E#),
      422 => to_slv(opcode_type, 16#05#),
      423 => to_slv(opcode_type, 16#11#),
      424 => to_slv(opcode_type, 16#09#),
      425 => to_slv(opcode_type, 16#0A#),
      426 => to_slv(opcode_type, 16#11#),
      427 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#07#),
      449 => to_slv(opcode_type, 16#08#),
      450 => to_slv(opcode_type, 16#03#),
      451 => to_slv(opcode_type, 16#07#),
      452 => to_slv(opcode_type, 16#10#),
      453 => to_slv(opcode_type, 16#11#),
      454 => to_slv(opcode_type, 16#02#),
      455 => to_slv(opcode_type, 16#06#),
      456 => to_slv(opcode_type, 16#0A#),
      457 => to_slv(opcode_type, 16#0E#),
      458 => to_slv(opcode_type, 16#0F#),
      459 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#04#),
      481 => to_slv(opcode_type, 16#08#),
      482 => to_slv(opcode_type, 16#03#),
      483 => to_slv(opcode_type, 16#09#),
      484 => to_slv(opcode_type, 16#0B#),
      485 => to_slv(opcode_type, 16#68#),
      486 => to_slv(opcode_type, 16#08#),
      487 => to_slv(opcode_type, 16#05#),
      488 => to_slv(opcode_type, 16#0B#),
      489 => to_slv(opcode_type, 16#05#),
      490 => to_slv(opcode_type, 16#0B#),
      491 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#06#),
      513 => to_slv(opcode_type, 16#05#),
      514 => to_slv(opcode_type, 16#01#),
      515 => to_slv(opcode_type, 16#05#),
      516 => to_slv(opcode_type, 16#11#),
      517 => to_slv(opcode_type, 16#01#),
      518 => to_slv(opcode_type, 16#07#),
      519 => to_slv(opcode_type, 16#04#),
      520 => to_slv(opcode_type, 16#0A#),
      521 => to_slv(opcode_type, 16#01#),
      522 => to_slv(opcode_type, 16#EE#),
      523 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#02#),
      545 => to_slv(opcode_type, 16#07#),
      546 => to_slv(opcode_type, 16#03#),
      547 => to_slv(opcode_type, 16#02#),
      548 => to_slv(opcode_type, 16#0F#),
      549 => to_slv(opcode_type, 16#06#),
      550 => to_slv(opcode_type, 16#04#),
      551 => to_slv(opcode_type, 16#0A#),
      552 => to_slv(opcode_type, 16#07#),
      553 => to_slv(opcode_type, 16#0C#),
      554 => to_slv(opcode_type, 16#0A#),
      555 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#02#),
      577 => to_slv(opcode_type, 16#07#),
      578 => to_slv(opcode_type, 16#09#),
      579 => to_slv(opcode_type, 16#05#),
      580 => to_slv(opcode_type, 16#B2#),
      581 => to_slv(opcode_type, 16#07#),
      582 => to_slv(opcode_type, 16#10#),
      583 => to_slv(opcode_type, 16#0C#),
      584 => to_slv(opcode_type, 16#09#),
      585 => to_slv(opcode_type, 16#0E#),
      586 => to_slv(opcode_type, 16#0C#),
      587 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#08#),
      609 => to_slv(opcode_type, 16#09#),
      610 => to_slv(opcode_type, 16#03#),
      611 => to_slv(opcode_type, 16#03#),
      612 => to_slv(opcode_type, 16#0C#),
      613 => to_slv(opcode_type, 16#04#),
      614 => to_slv(opcode_type, 16#02#),
      615 => to_slv(opcode_type, 16#11#),
      616 => to_slv(opcode_type, 16#06#),
      617 => to_slv(opcode_type, 16#0B#),
      618 => to_slv(opcode_type, 16#0D#),
      619 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#03#),
      641 => to_slv(opcode_type, 16#07#),
      642 => to_slv(opcode_type, 16#07#),
      643 => to_slv(opcode_type, 16#05#),
      644 => to_slv(opcode_type, 16#0F#),
      645 => to_slv(opcode_type, 16#07#),
      646 => to_slv(opcode_type, 16#0B#),
      647 => to_slv(opcode_type, 16#0D#),
      648 => to_slv(opcode_type, 16#08#),
      649 => to_slv(opcode_type, 16#10#),
      650 => to_slv(opcode_type, 16#0E#),
      651 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#03#),
      673 => to_slv(opcode_type, 16#08#),
      674 => to_slv(opcode_type, 16#08#),
      675 => to_slv(opcode_type, 16#02#),
      676 => to_slv(opcode_type, 16#69#),
      677 => to_slv(opcode_type, 16#04#),
      678 => to_slv(opcode_type, 16#30#),
      679 => to_slv(opcode_type, 16#06#),
      680 => to_slv(opcode_type, 16#03#),
      681 => to_slv(opcode_type, 16#0E#),
      682 => to_slv(opcode_type, 16#10#),
      683 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#04#),
      705 => to_slv(opcode_type, 16#08#),
      706 => to_slv(opcode_type, 16#02#),
      707 => to_slv(opcode_type, 16#05#),
      708 => to_slv(opcode_type, 16#0B#),
      709 => to_slv(opcode_type, 16#07#),
      710 => to_slv(opcode_type, 16#08#),
      711 => to_slv(opcode_type, 16#0F#),
      712 => to_slv(opcode_type, 16#E7#),
      713 => to_slv(opcode_type, 16#01#),
      714 => to_slv(opcode_type, 16#C0#),
      715 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#06#),
      737 => to_slv(opcode_type, 16#06#),
      738 => to_slv(opcode_type, 16#05#),
      739 => to_slv(opcode_type, 16#08#),
      740 => to_slv(opcode_type, 16#10#),
      741 => to_slv(opcode_type, 16#0A#),
      742 => to_slv(opcode_type, 16#09#),
      743 => to_slv(opcode_type, 16#04#),
      744 => to_slv(opcode_type, 16#11#),
      745 => to_slv(opcode_type, 16#F4#),
      746 => to_slv(opcode_type, 16#10#),
      747 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#04#),
      769 => to_slv(opcode_type, 16#06#),
      770 => to_slv(opcode_type, 16#01#),
      771 => to_slv(opcode_type, 16#05#),
      772 => to_slv(opcode_type, 16#0A#),
      773 => to_slv(opcode_type, 16#06#),
      774 => to_slv(opcode_type, 16#09#),
      775 => to_slv(opcode_type, 16#0B#),
      776 => to_slv(opcode_type, 16#0D#),
      777 => to_slv(opcode_type, 16#01#),
      778 => to_slv(opcode_type, 16#11#),
      779 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#07#),
      801 => to_slv(opcode_type, 16#09#),
      802 => to_slv(opcode_type, 16#04#),
      803 => to_slv(opcode_type, 16#03#),
      804 => to_slv(opcode_type, 16#3A#),
      805 => to_slv(opcode_type, 16#09#),
      806 => to_slv(opcode_type, 16#05#),
      807 => to_slv(opcode_type, 16#0A#),
      808 => to_slv(opcode_type, 16#03#),
      809 => to_slv(opcode_type, 16#0B#),
      810 => to_slv(opcode_type, 16#0B#),
      811 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#04#),
      833 => to_slv(opcode_type, 16#08#),
      834 => to_slv(opcode_type, 16#09#),
      835 => to_slv(opcode_type, 16#08#),
      836 => to_slv(opcode_type, 16#0B#),
      837 => to_slv(opcode_type, 16#0B#),
      838 => to_slv(opcode_type, 16#06#),
      839 => to_slv(opcode_type, 16#10#),
      840 => to_slv(opcode_type, 16#10#),
      841 => to_slv(opcode_type, 16#05#),
      842 => to_slv(opcode_type, 16#0C#),
      843 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#02#),
      865 => to_slv(opcode_type, 16#08#),
      866 => to_slv(opcode_type, 16#01#),
      867 => to_slv(opcode_type, 16#01#),
      868 => to_slv(opcode_type, 16#0C#),
      869 => to_slv(opcode_type, 16#09#),
      870 => to_slv(opcode_type, 16#03#),
      871 => to_slv(opcode_type, 16#0F#),
      872 => to_slv(opcode_type, 16#09#),
      873 => to_slv(opcode_type, 16#10#),
      874 => to_slv(opcode_type, 16#0E#),
      875 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#02#),
      898 => to_slv(opcode_type, 16#05#),
      899 => to_slv(opcode_type, 16#07#),
      900 => to_slv(opcode_type, 16#0A#),
      901 => to_slv(opcode_type, 16#0E#),
      902 => to_slv(opcode_type, 16#02#),
      903 => to_slv(opcode_type, 16#04#),
      904 => to_slv(opcode_type, 16#09#),
      905 => to_slv(opcode_type, 16#0C#),
      906 => to_slv(opcode_type, 16#0C#),
      907 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#04#),
      929 => to_slv(opcode_type, 16#08#),
      930 => to_slv(opcode_type, 16#05#),
      931 => to_slv(opcode_type, 16#01#),
      932 => to_slv(opcode_type, 16#0A#),
      933 => to_slv(opcode_type, 16#06#),
      934 => to_slv(opcode_type, 16#06#),
      935 => to_slv(opcode_type, 16#11#),
      936 => to_slv(opcode_type, 16#0A#),
      937 => to_slv(opcode_type, 16#02#),
      938 => to_slv(opcode_type, 16#0C#),
      939 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#05#),
      961 => to_slv(opcode_type, 16#07#),
      962 => to_slv(opcode_type, 16#05#),
      963 => to_slv(opcode_type, 16#04#),
      964 => to_slv(opcode_type, 16#0A#),
      965 => to_slv(opcode_type, 16#06#),
      966 => to_slv(opcode_type, 16#02#),
      967 => to_slv(opcode_type, 16#0B#),
      968 => to_slv(opcode_type, 16#09#),
      969 => to_slv(opcode_type, 16#11#),
      970 => to_slv(opcode_type, 16#0B#),
      971 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#05#),
      993 => to_slv(opcode_type, 16#06#),
      994 => to_slv(opcode_type, 16#03#),
      995 => to_slv(opcode_type, 16#09#),
      996 => to_slv(opcode_type, 16#11#),
      997 => to_slv(opcode_type, 16#0E#),
      998 => to_slv(opcode_type, 16#08#),
      999 => to_slv(opcode_type, 16#09#),
      1000 => to_slv(opcode_type, 16#7F#),
      1001 => to_slv(opcode_type, 16#B1#),
      1002 => to_slv(opcode_type, 16#0B#),
      1003 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#03#),
      1025 => to_slv(opcode_type, 16#08#),
      1026 => to_slv(opcode_type, 16#08#),
      1027 => to_slv(opcode_type, 16#06#),
      1028 => to_slv(opcode_type, 16#10#),
      1029 => to_slv(opcode_type, 16#63#),
      1030 => to_slv(opcode_type, 16#02#),
      1031 => to_slv(opcode_type, 16#0D#),
      1032 => to_slv(opcode_type, 16#02#),
      1033 => to_slv(opcode_type, 16#01#),
      1034 => to_slv(opcode_type, 16#0B#),
      1035 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#01#),
      1057 => to_slv(opcode_type, 16#07#),
      1058 => to_slv(opcode_type, 16#03#),
      1059 => to_slv(opcode_type, 16#07#),
      1060 => to_slv(opcode_type, 16#0E#),
      1061 => to_slv(opcode_type, 16#0A#),
      1062 => to_slv(opcode_type, 16#07#),
      1063 => to_slv(opcode_type, 16#01#),
      1064 => to_slv(opcode_type, 16#11#),
      1065 => to_slv(opcode_type, 16#01#),
      1066 => to_slv(opcode_type, 16#0B#),
      1067 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#08#),
      1089 => to_slv(opcode_type, 16#02#),
      1090 => to_slv(opcode_type, 16#04#),
      1091 => to_slv(opcode_type, 16#09#),
      1092 => to_slv(opcode_type, 16#0B#),
      1093 => to_slv(opcode_type, 16#0C#),
      1094 => to_slv(opcode_type, 16#01#),
      1095 => to_slv(opcode_type, 16#07#),
      1096 => to_slv(opcode_type, 16#02#),
      1097 => to_slv(opcode_type, 16#0D#),
      1098 => to_slv(opcode_type, 16#0A#),
      1099 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#09#),
      1121 => to_slv(opcode_type, 16#02#),
      1122 => to_slv(opcode_type, 16#08#),
      1123 => to_slv(opcode_type, 16#02#),
      1124 => to_slv(opcode_type, 16#0C#),
      1125 => to_slv(opcode_type, 16#07#),
      1126 => to_slv(opcode_type, 16#0B#),
      1127 => to_slv(opcode_type, 16#10#),
      1128 => to_slv(opcode_type, 16#07#),
      1129 => to_slv(opcode_type, 16#0B#),
      1130 => to_slv(opcode_type, 16#0F#),
      1131 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#03#),
      1153 => to_slv(opcode_type, 16#07#),
      1154 => to_slv(opcode_type, 16#05#),
      1155 => to_slv(opcode_type, 16#07#),
      1156 => to_slv(opcode_type, 16#0F#),
      1157 => to_slv(opcode_type, 16#0F#),
      1158 => to_slv(opcode_type, 16#08#),
      1159 => to_slv(opcode_type, 16#03#),
      1160 => to_slv(opcode_type, 16#10#),
      1161 => to_slv(opcode_type, 16#04#),
      1162 => to_slv(opcode_type, 16#0E#),
      1163 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#03#),
      1185 => to_slv(opcode_type, 16#06#),
      1186 => to_slv(opcode_type, 16#03#),
      1187 => to_slv(opcode_type, 16#08#),
      1188 => to_slv(opcode_type, 16#0E#),
      1189 => to_slv(opcode_type, 16#0E#),
      1190 => to_slv(opcode_type, 16#06#),
      1191 => to_slv(opcode_type, 16#06#),
      1192 => to_slv(opcode_type, 16#11#),
      1193 => to_slv(opcode_type, 16#0B#),
      1194 => to_slv(opcode_type, 16#0F#),
      1195 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#05#),
      1217 => to_slv(opcode_type, 16#06#),
      1218 => to_slv(opcode_type, 16#08#),
      1219 => to_slv(opcode_type, 16#07#),
      1220 => to_slv(opcode_type, 16#F1#),
      1221 => to_slv(opcode_type, 16#0C#),
      1222 => to_slv(opcode_type, 16#03#),
      1223 => to_slv(opcode_type, 16#0A#),
      1224 => to_slv(opcode_type, 16#06#),
      1225 => to_slv(opcode_type, 16#0D#),
      1226 => to_slv(opcode_type, 16#0F#),
      1227 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#04#),
      1249 => to_slv(opcode_type, 16#08#),
      1250 => to_slv(opcode_type, 16#03#),
      1251 => to_slv(opcode_type, 16#06#),
      1252 => to_slv(opcode_type, 16#0E#),
      1253 => to_slv(opcode_type, 16#0C#),
      1254 => to_slv(opcode_type, 16#09#),
      1255 => to_slv(opcode_type, 16#03#),
      1256 => to_slv(opcode_type, 16#0B#),
      1257 => to_slv(opcode_type, 16#01#),
      1258 => to_slv(opcode_type, 16#0C#),
      1259 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#07#),
      1281 => to_slv(opcode_type, 16#01#),
      1282 => to_slv(opcode_type, 16#09#),
      1283 => to_slv(opcode_type, 16#08#),
      1284 => to_slv(opcode_type, 16#0A#),
      1285 => to_slv(opcode_type, 16#0D#),
      1286 => to_slv(opcode_type, 16#02#),
      1287 => to_slv(opcode_type, 16#0E#),
      1288 => to_slv(opcode_type, 16#01#),
      1289 => to_slv(opcode_type, 16#01#),
      1290 => to_slv(opcode_type, 16#0F#),
      1291 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#05#),
      1313 => to_slv(opcode_type, 16#09#),
      1314 => to_slv(opcode_type, 16#08#),
      1315 => to_slv(opcode_type, 16#03#),
      1316 => to_slv(opcode_type, 16#11#),
      1317 => to_slv(opcode_type, 16#07#),
      1318 => to_slv(opcode_type, 16#11#),
      1319 => to_slv(opcode_type, 16#0C#),
      1320 => to_slv(opcode_type, 16#08#),
      1321 => to_slv(opcode_type, 16#0C#),
      1322 => to_slv(opcode_type, 16#0D#),
      1323 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#02#),
      1345 => to_slv(opcode_type, 16#06#),
      1346 => to_slv(opcode_type, 16#02#),
      1347 => to_slv(opcode_type, 16#02#),
      1348 => to_slv(opcode_type, 16#0A#),
      1349 => to_slv(opcode_type, 16#09#),
      1350 => to_slv(opcode_type, 16#03#),
      1351 => to_slv(opcode_type, 16#12#),
      1352 => to_slv(opcode_type, 16#06#),
      1353 => to_slv(opcode_type, 16#49#),
      1354 => to_slv(opcode_type, 16#0D#),
      1355 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#08#),
      1377 => to_slv(opcode_type, 16#06#),
      1378 => to_slv(opcode_type, 16#07#),
      1379 => to_slv(opcode_type, 16#05#),
      1380 => to_slv(opcode_type, 16#0C#),
      1381 => to_slv(opcode_type, 16#01#),
      1382 => to_slv(opcode_type, 16#0A#),
      1383 => to_slv(opcode_type, 16#06#),
      1384 => to_slv(opcode_type, 16#10#),
      1385 => to_slv(opcode_type, 16#0A#),
      1386 => to_slv(opcode_type, 16#0B#),
      1387 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#07#),
      1409 => to_slv(opcode_type, 16#03#),
      1410 => to_slv(opcode_type, 16#06#),
      1411 => to_slv(opcode_type, 16#08#),
      1412 => to_slv(opcode_type, 16#0E#),
      1413 => to_slv(opcode_type, 16#0F#),
      1414 => to_slv(opcode_type, 16#09#),
      1415 => to_slv(opcode_type, 16#0B#),
      1416 => to_slv(opcode_type, 16#D3#),
      1417 => to_slv(opcode_type, 16#04#),
      1418 => to_slv(opcode_type, 16#0C#),
      1419 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#06#),
      1441 => to_slv(opcode_type, 16#07#),
      1442 => to_slv(opcode_type, 16#01#),
      1443 => to_slv(opcode_type, 16#08#),
      1444 => to_slv(opcode_type, 16#11#),
      1445 => to_slv(opcode_type, 16#0F#),
      1446 => to_slv(opcode_type, 16#05#),
      1447 => to_slv(opcode_type, 16#09#),
      1448 => to_slv(opcode_type, 16#0F#),
      1449 => to_slv(opcode_type, 16#0C#),
      1450 => to_slv(opcode_type, 16#11#),
      1451 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#05#),
      1473 => to_slv(opcode_type, 16#08#),
      1474 => to_slv(opcode_type, 16#04#),
      1475 => to_slv(opcode_type, 16#01#),
      1476 => to_slv(opcode_type, 16#0D#),
      1477 => to_slv(opcode_type, 16#06#),
      1478 => to_slv(opcode_type, 16#03#),
      1479 => to_slv(opcode_type, 16#11#),
      1480 => to_slv(opcode_type, 16#08#),
      1481 => to_slv(opcode_type, 16#0B#),
      1482 => to_slv(opcode_type, 16#0E#),
      1483 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#01#),
      1505 => to_slv(opcode_type, 16#08#),
      1506 => to_slv(opcode_type, 16#04#),
      1507 => to_slv(opcode_type, 16#04#),
      1508 => to_slv(opcode_type, 16#11#),
      1509 => to_slv(opcode_type, 16#09#),
      1510 => to_slv(opcode_type, 16#06#),
      1511 => to_slv(opcode_type, 16#0E#),
      1512 => to_slv(opcode_type, 16#0B#),
      1513 => to_slv(opcode_type, 16#01#),
      1514 => to_slv(opcode_type, 16#0C#),
      1515 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#03#),
      1537 => to_slv(opcode_type, 16#06#),
      1538 => to_slv(opcode_type, 16#08#),
      1539 => to_slv(opcode_type, 16#09#),
      1540 => to_slv(opcode_type, 16#0A#),
      1541 => to_slv(opcode_type, 16#0A#),
      1542 => to_slv(opcode_type, 16#09#),
      1543 => to_slv(opcode_type, 16#83#),
      1544 => to_slv(opcode_type, 16#0A#),
      1545 => to_slv(opcode_type, 16#05#),
      1546 => to_slv(opcode_type, 16#0C#),
      1547 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#04#),
      1569 => to_slv(opcode_type, 16#08#),
      1570 => to_slv(opcode_type, 16#07#),
      1571 => to_slv(opcode_type, 16#01#),
      1572 => to_slv(opcode_type, 16#0C#),
      1573 => to_slv(opcode_type, 16#07#),
      1574 => to_slv(opcode_type, 16#0E#),
      1575 => to_slv(opcode_type, 16#0C#),
      1576 => to_slv(opcode_type, 16#06#),
      1577 => to_slv(opcode_type, 16#10#),
      1578 => to_slv(opcode_type, 16#0C#),
      1579 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#04#),
      1601 => to_slv(opcode_type, 16#09#),
      1602 => to_slv(opcode_type, 16#06#),
      1603 => to_slv(opcode_type, 16#01#),
      1604 => to_slv(opcode_type, 16#0C#),
      1605 => to_slv(opcode_type, 16#02#),
      1606 => to_slv(opcode_type, 16#11#),
      1607 => to_slv(opcode_type, 16#04#),
      1608 => to_slv(opcode_type, 16#09#),
      1609 => to_slv(opcode_type, 16#0F#),
      1610 => to_slv(opcode_type, 16#6D#),
      1611 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#06#),
      1633 => to_slv(opcode_type, 16#06#),
      1634 => to_slv(opcode_type, 16#04#),
      1635 => to_slv(opcode_type, 16#03#),
      1636 => to_slv(opcode_type, 16#0D#),
      1637 => to_slv(opcode_type, 16#09#),
      1638 => to_slv(opcode_type, 16#04#),
      1639 => to_slv(opcode_type, 16#11#),
      1640 => to_slv(opcode_type, 16#05#),
      1641 => to_slv(opcode_type, 16#0B#),
      1642 => to_slv(opcode_type, 16#10#),
      1643 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#08#),
      1666 => to_slv(opcode_type, 16#02#),
      1667 => to_slv(opcode_type, 16#03#),
      1668 => to_slv(opcode_type, 16#10#),
      1669 => to_slv(opcode_type, 16#05#),
      1670 => to_slv(opcode_type, 16#09#),
      1671 => to_slv(opcode_type, 16#10#),
      1672 => to_slv(opcode_type, 16#0D#),
      1673 => to_slv(opcode_type, 16#05#),
      1674 => to_slv(opcode_type, 16#0B#),
      1675 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#05#),
      1697 => to_slv(opcode_type, 16#07#),
      1698 => to_slv(opcode_type, 16#08#),
      1699 => to_slv(opcode_type, 16#05#),
      1700 => to_slv(opcode_type, 16#0F#),
      1701 => to_slv(opcode_type, 16#02#),
      1702 => to_slv(opcode_type, 16#0D#),
      1703 => to_slv(opcode_type, 16#08#),
      1704 => to_slv(opcode_type, 16#05#),
      1705 => to_slv(opcode_type, 16#0A#),
      1706 => to_slv(opcode_type, 16#0B#),
      1707 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#05#),
      1729 => to_slv(opcode_type, 16#07#),
      1730 => to_slv(opcode_type, 16#06#),
      1731 => to_slv(opcode_type, 16#02#),
      1732 => to_slv(opcode_type, 16#0B#),
      1733 => to_slv(opcode_type, 16#04#),
      1734 => to_slv(opcode_type, 16#0A#),
      1735 => to_slv(opcode_type, 16#07#),
      1736 => to_slv(opcode_type, 16#01#),
      1737 => to_slv(opcode_type, 16#11#),
      1738 => to_slv(opcode_type, 16#0B#),
      1739 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#04#),
      1761 => to_slv(opcode_type, 16#09#),
      1762 => to_slv(opcode_type, 16#09#),
      1763 => to_slv(opcode_type, 16#05#),
      1764 => to_slv(opcode_type, 16#11#),
      1765 => to_slv(opcode_type, 16#09#),
      1766 => to_slv(opcode_type, 16#11#),
      1767 => to_slv(opcode_type, 16#0E#),
      1768 => to_slv(opcode_type, 16#04#),
      1769 => to_slv(opcode_type, 16#01#),
      1770 => to_slv(opcode_type, 16#0F#),
      1771 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#05#),
      1793 => to_slv(opcode_type, 16#07#),
      1794 => to_slv(opcode_type, 16#03#),
      1795 => to_slv(opcode_type, 16#04#),
      1796 => to_slv(opcode_type, 16#10#),
      1797 => to_slv(opcode_type, 16#07#),
      1798 => to_slv(opcode_type, 16#03#),
      1799 => to_slv(opcode_type, 16#0A#),
      1800 => to_slv(opcode_type, 16#08#),
      1801 => to_slv(opcode_type, 16#0D#),
      1802 => to_slv(opcode_type, 16#0E#),
      1803 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#07#),
      1825 => to_slv(opcode_type, 16#02#),
      1826 => to_slv(opcode_type, 16#04#),
      1827 => to_slv(opcode_type, 16#03#),
      1828 => to_slv(opcode_type, 16#0E#),
      1829 => to_slv(opcode_type, 16#02#),
      1830 => to_slv(opcode_type, 16#06#),
      1831 => to_slv(opcode_type, 16#07#),
      1832 => to_slv(opcode_type, 16#33#),
      1833 => to_slv(opcode_type, 16#0F#),
      1834 => to_slv(opcode_type, 16#0A#),
      1835 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#03#),
      1857 => to_slv(opcode_type, 16#08#),
      1858 => to_slv(opcode_type, 16#09#),
      1859 => to_slv(opcode_type, 16#08#),
      1860 => to_slv(opcode_type, 16#DB#),
      1861 => to_slv(opcode_type, 16#10#),
      1862 => to_slv(opcode_type, 16#07#),
      1863 => to_slv(opcode_type, 16#0D#),
      1864 => to_slv(opcode_type, 16#10#),
      1865 => to_slv(opcode_type, 16#03#),
      1866 => to_slv(opcode_type, 16#10#),
      1867 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#03#),
      1889 => to_slv(opcode_type, 16#07#),
      1890 => to_slv(opcode_type, 16#09#),
      1891 => to_slv(opcode_type, 16#07#),
      1892 => to_slv(opcode_type, 16#0F#),
      1893 => to_slv(opcode_type, 16#0C#),
      1894 => to_slv(opcode_type, 16#03#),
      1895 => to_slv(opcode_type, 16#0C#),
      1896 => to_slv(opcode_type, 16#06#),
      1897 => to_slv(opcode_type, 16#0D#),
      1898 => to_slv(opcode_type, 16#0F#),
      1899 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#02#),
      1921 => to_slv(opcode_type, 16#08#),
      1922 => to_slv(opcode_type, 16#04#),
      1923 => to_slv(opcode_type, 16#03#),
      1924 => to_slv(opcode_type, 16#11#),
      1925 => to_slv(opcode_type, 16#08#),
      1926 => to_slv(opcode_type, 16#04#),
      1927 => to_slv(opcode_type, 16#0E#),
      1928 => to_slv(opcode_type, 16#09#),
      1929 => to_slv(opcode_type, 16#0A#),
      1930 => to_slv(opcode_type, 16#11#),
      1931 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#08#),
      1953 => to_slv(opcode_type, 16#03#),
      1954 => to_slv(opcode_type, 16#01#),
      1955 => to_slv(opcode_type, 16#05#),
      1956 => to_slv(opcode_type, 16#0D#),
      1957 => to_slv(opcode_type, 16#02#),
      1958 => to_slv(opcode_type, 16#07#),
      1959 => to_slv(opcode_type, 16#07#),
      1960 => to_slv(opcode_type, 16#0F#),
      1961 => to_slv(opcode_type, 16#11#),
      1962 => to_slv(opcode_type, 16#0D#),
      1963 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#03#),
      1985 => to_slv(opcode_type, 16#09#),
      1986 => to_slv(opcode_type, 16#01#),
      1987 => to_slv(opcode_type, 16#07#),
      1988 => to_slv(opcode_type, 16#0B#),
      1989 => to_slv(opcode_type, 16#0E#),
      1990 => to_slv(opcode_type, 16#09#),
      1991 => to_slv(opcode_type, 16#03#),
      1992 => to_slv(opcode_type, 16#0A#),
      1993 => to_slv(opcode_type, 16#02#),
      1994 => to_slv(opcode_type, 16#0A#),
      1995 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#08#),
      2017 => to_slv(opcode_type, 16#05#),
      2018 => to_slv(opcode_type, 16#03#),
      2019 => to_slv(opcode_type, 16#04#),
      2020 => to_slv(opcode_type, 16#0D#),
      2021 => to_slv(opcode_type, 16#04#),
      2022 => to_slv(opcode_type, 16#09#),
      2023 => to_slv(opcode_type, 16#03#),
      2024 => to_slv(opcode_type, 16#11#),
      2025 => to_slv(opcode_type, 16#01#),
      2026 => to_slv(opcode_type, 16#0A#),
      2027 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#08#),
      2049 => to_slv(opcode_type, 16#03#),
      2050 => to_slv(opcode_type, 16#09#),
      2051 => to_slv(opcode_type, 16#09#),
      2052 => to_slv(opcode_type, 16#10#),
      2053 => to_slv(opcode_type, 16#0B#),
      2054 => to_slv(opcode_type, 16#09#),
      2055 => to_slv(opcode_type, 16#0A#),
      2056 => to_slv(opcode_type, 16#10#),
      2057 => to_slv(opcode_type, 16#05#),
      2058 => to_slv(opcode_type, 16#0A#),
      2059 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#06#),
      2081 => to_slv(opcode_type, 16#07#),
      2082 => to_slv(opcode_type, 16#01#),
      2083 => to_slv(opcode_type, 16#09#),
      2084 => to_slv(opcode_type, 16#C8#),
      2085 => to_slv(opcode_type, 16#0F#),
      2086 => to_slv(opcode_type, 16#08#),
      2087 => to_slv(opcode_type, 16#04#),
      2088 => to_slv(opcode_type, 16#0A#),
      2089 => to_slv(opcode_type, 16#0C#),
      2090 => to_slv(opcode_type, 16#0B#),
      2091 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#05#),
      2113 => to_slv(opcode_type, 16#09#),
      2114 => to_slv(opcode_type, 16#05#),
      2115 => to_slv(opcode_type, 16#03#),
      2116 => to_slv(opcode_type, 16#11#),
      2117 => to_slv(opcode_type, 16#08#),
      2118 => to_slv(opcode_type, 16#05#),
      2119 => to_slv(opcode_type, 16#10#),
      2120 => to_slv(opcode_type, 16#08#),
      2121 => to_slv(opcode_type, 16#61#),
      2122 => to_slv(opcode_type, 16#10#),
      2123 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#03#),
      2145 => to_slv(opcode_type, 16#09#),
      2146 => to_slv(opcode_type, 16#08#),
      2147 => to_slv(opcode_type, 16#09#),
      2148 => to_slv(opcode_type, 16#0A#),
      2149 => to_slv(opcode_type, 16#11#),
      2150 => to_slv(opcode_type, 16#04#),
      2151 => to_slv(opcode_type, 16#0B#),
      2152 => to_slv(opcode_type, 16#01#),
      2153 => to_slv(opcode_type, 16#05#),
      2154 => to_slv(opcode_type, 16#69#),
      2155 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#01#),
      2177 => to_slv(opcode_type, 16#07#),
      2178 => to_slv(opcode_type, 16#01#),
      2179 => to_slv(opcode_type, 16#05#),
      2180 => to_slv(opcode_type, 16#10#),
      2181 => to_slv(opcode_type, 16#08#),
      2182 => to_slv(opcode_type, 16#09#),
      2183 => to_slv(opcode_type, 16#0A#),
      2184 => to_slv(opcode_type, 16#A0#),
      2185 => to_slv(opcode_type, 16#02#),
      2186 => to_slv(opcode_type, 16#0E#),
      2187 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#09#),
      2209 => to_slv(opcode_type, 16#01#),
      2210 => to_slv(opcode_type, 16#01#),
      2211 => to_slv(opcode_type, 16#03#),
      2212 => to_slv(opcode_type, 16#10#),
      2213 => to_slv(opcode_type, 16#03#),
      2214 => to_slv(opcode_type, 16#08#),
      2215 => to_slv(opcode_type, 16#05#),
      2216 => to_slv(opcode_type, 16#10#),
      2217 => to_slv(opcode_type, 16#03#),
      2218 => to_slv(opcode_type, 16#0A#),
      2219 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#08#),
      2241 => to_slv(opcode_type, 16#09#),
      2242 => to_slv(opcode_type, 16#04#),
      2243 => to_slv(opcode_type, 16#06#),
      2244 => to_slv(opcode_type, 16#0D#),
      2245 => to_slv(opcode_type, 16#6F#),
      2246 => to_slv(opcode_type, 16#09#),
      2247 => to_slv(opcode_type, 16#02#),
      2248 => to_slv(opcode_type, 16#0B#),
      2249 => to_slv(opcode_type, 16#0D#),
      2250 => to_slv(opcode_type, 16#0E#),
      2251 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#04#),
      2273 => to_slv(opcode_type, 16#09#),
      2274 => to_slv(opcode_type, 16#05#),
      2275 => to_slv(opcode_type, 16#08#),
      2276 => to_slv(opcode_type, 16#0F#),
      2277 => to_slv(opcode_type, 16#11#),
      2278 => to_slv(opcode_type, 16#06#),
      2279 => to_slv(opcode_type, 16#03#),
      2280 => to_slv(opcode_type, 16#11#),
      2281 => to_slv(opcode_type, 16#02#),
      2282 => to_slv(opcode_type, 16#0B#),
      2283 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#05#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#01#),
      2307 => to_slv(opcode_type, 16#02#),
      2308 => to_slv(opcode_type, 16#0D#),
      2309 => to_slv(opcode_type, 16#08#),
      2310 => to_slv(opcode_type, 16#03#),
      2311 => to_slv(opcode_type, 16#0E#),
      2312 => to_slv(opcode_type, 16#06#),
      2313 => to_slv(opcode_type, 16#11#),
      2314 => to_slv(opcode_type, 16#11#),
      2315 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#08#),
      2337 => to_slv(opcode_type, 16#06#),
      2338 => to_slv(opcode_type, 16#08#),
      2339 => to_slv(opcode_type, 16#07#),
      2340 => to_slv(opcode_type, 16#11#),
      2341 => to_slv(opcode_type, 16#0C#),
      2342 => to_slv(opcode_type, 16#04#),
      2343 => to_slv(opcode_type, 16#0D#),
      2344 => to_slv(opcode_type, 16#05#),
      2345 => to_slv(opcode_type, 16#0B#),
      2346 => to_slv(opcode_type, 16#10#),
      2347 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#06#),
      2369 => to_slv(opcode_type, 16#03#),
      2370 => to_slv(opcode_type, 16#09#),
      2371 => to_slv(opcode_type, 16#03#),
      2372 => to_slv(opcode_type, 16#10#),
      2373 => to_slv(opcode_type, 16#07#),
      2374 => to_slv(opcode_type, 16#0A#),
      2375 => to_slv(opcode_type, 16#0B#),
      2376 => to_slv(opcode_type, 16#09#),
      2377 => to_slv(opcode_type, 16#10#),
      2378 => to_slv(opcode_type, 16#13#),
      2379 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#07#),
      2401 => to_slv(opcode_type, 16#02#),
      2402 => to_slv(opcode_type, 16#02#),
      2403 => to_slv(opcode_type, 16#02#),
      2404 => to_slv(opcode_type, 16#0B#),
      2405 => to_slv(opcode_type, 16#07#),
      2406 => to_slv(opcode_type, 16#02#),
      2407 => to_slv(opcode_type, 16#06#),
      2408 => to_slv(opcode_type, 16#0A#),
      2409 => to_slv(opcode_type, 16#0B#),
      2410 => to_slv(opcode_type, 16#0E#),
      2411 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#06#),
      2433 => to_slv(opcode_type, 16#08#),
      2434 => to_slv(opcode_type, 16#05#),
      2435 => to_slv(opcode_type, 16#05#),
      2436 => to_slv(opcode_type, 16#89#),
      2437 => to_slv(opcode_type, 16#06#),
      2438 => to_slv(opcode_type, 16#01#),
      2439 => to_slv(opcode_type, 16#0E#),
      2440 => to_slv(opcode_type, 16#01#),
      2441 => to_slv(opcode_type, 16#D5#),
      2442 => to_slv(opcode_type, 16#0F#),
      2443 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#03#),
      2465 => to_slv(opcode_type, 16#09#),
      2466 => to_slv(opcode_type, 16#08#),
      2467 => to_slv(opcode_type, 16#09#),
      2468 => to_slv(opcode_type, 16#0D#),
      2469 => to_slv(opcode_type, 16#0A#),
      2470 => to_slv(opcode_type, 16#03#),
      2471 => to_slv(opcode_type, 16#10#),
      2472 => to_slv(opcode_type, 16#02#),
      2473 => to_slv(opcode_type, 16#05#),
      2474 => to_slv(opcode_type, 16#0D#),
      2475 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#01#),
      2497 => to_slv(opcode_type, 16#09#),
      2498 => to_slv(opcode_type, 16#01#),
      2499 => to_slv(opcode_type, 16#07#),
      2500 => to_slv(opcode_type, 16#0B#),
      2501 => to_slv(opcode_type, 16#0A#),
      2502 => to_slv(opcode_type, 16#08#),
      2503 => to_slv(opcode_type, 16#01#),
      2504 => to_slv(opcode_type, 16#11#),
      2505 => to_slv(opcode_type, 16#01#),
      2506 => to_slv(opcode_type, 16#EB#),
      2507 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#01#),
      2529 => to_slv(opcode_type, 16#06#),
      2530 => to_slv(opcode_type, 16#02#),
      2531 => to_slv(opcode_type, 16#08#),
      2532 => to_slv(opcode_type, 16#99#),
      2533 => to_slv(opcode_type, 16#11#),
      2534 => to_slv(opcode_type, 16#07#),
      2535 => to_slv(opcode_type, 16#09#),
      2536 => to_slv(opcode_type, 16#0C#),
      2537 => to_slv(opcode_type, 16#0B#),
      2538 => to_slv(opcode_type, 16#0B#),
      2539 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#02#),
      2561 => to_slv(opcode_type, 16#08#),
      2562 => to_slv(opcode_type, 16#04#),
      2563 => to_slv(opcode_type, 16#07#),
      2564 => to_slv(opcode_type, 16#0B#),
      2565 => to_slv(opcode_type, 16#0F#),
      2566 => to_slv(opcode_type, 16#08#),
      2567 => to_slv(opcode_type, 16#07#),
      2568 => to_slv(opcode_type, 16#0E#),
      2569 => to_slv(opcode_type, 16#11#),
      2570 => to_slv(opcode_type, 16#0E#),
      2571 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#02#),
      2593 => to_slv(opcode_type, 16#07#),
      2594 => to_slv(opcode_type, 16#01#),
      2595 => to_slv(opcode_type, 16#02#),
      2596 => to_slv(opcode_type, 16#0E#),
      2597 => to_slv(opcode_type, 16#09#),
      2598 => to_slv(opcode_type, 16#09#),
      2599 => to_slv(opcode_type, 16#11#),
      2600 => to_slv(opcode_type, 16#9B#),
      2601 => to_slv(opcode_type, 16#04#),
      2602 => to_slv(opcode_type, 16#0C#),
      2603 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#05#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#04#),
      2627 => to_slv(opcode_type, 16#01#),
      2628 => to_slv(opcode_type, 16#0F#),
      2629 => to_slv(opcode_type, 16#06#),
      2630 => to_slv(opcode_type, 16#04#),
      2631 => to_slv(opcode_type, 16#0B#),
      2632 => to_slv(opcode_type, 16#06#),
      2633 => to_slv(opcode_type, 16#11#),
      2634 => to_slv(opcode_type, 16#10#),
      2635 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#04#),
      2657 => to_slv(opcode_type, 16#06#),
      2658 => to_slv(opcode_type, 16#08#),
      2659 => to_slv(opcode_type, 16#06#),
      2660 => to_slv(opcode_type, 16#0B#),
      2661 => to_slv(opcode_type, 16#11#),
      2662 => to_slv(opcode_type, 16#06#),
      2663 => to_slv(opcode_type, 16#0E#),
      2664 => to_slv(opcode_type, 16#0F#),
      2665 => to_slv(opcode_type, 16#01#),
      2666 => to_slv(opcode_type, 16#5D#),
      2667 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#02#),
      2689 => to_slv(opcode_type, 16#06#),
      2690 => to_slv(opcode_type, 16#01#),
      2691 => to_slv(opcode_type, 16#07#),
      2692 => to_slv(opcode_type, 16#10#),
      2693 => to_slv(opcode_type, 16#11#),
      2694 => to_slv(opcode_type, 16#06#),
      2695 => to_slv(opcode_type, 16#06#),
      2696 => to_slv(opcode_type, 16#0D#),
      2697 => to_slv(opcode_type, 16#0D#),
      2698 => to_slv(opcode_type, 16#0A#),
      2699 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#05#),
      2721 => to_slv(opcode_type, 16#07#),
      2722 => to_slv(opcode_type, 16#07#),
      2723 => to_slv(opcode_type, 16#04#),
      2724 => to_slv(opcode_type, 16#10#),
      2725 => to_slv(opcode_type, 16#03#),
      2726 => to_slv(opcode_type, 16#0C#),
      2727 => to_slv(opcode_type, 16#01#),
      2728 => to_slv(opcode_type, 16#08#),
      2729 => to_slv(opcode_type, 16#0A#),
      2730 => to_slv(opcode_type, 16#0B#),
      2731 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#07#),
      2753 => to_slv(opcode_type, 16#07#),
      2754 => to_slv(opcode_type, 16#04#),
      2755 => to_slv(opcode_type, 16#04#),
      2756 => to_slv(opcode_type, 16#0F#),
      2757 => to_slv(opcode_type, 16#09#),
      2758 => to_slv(opcode_type, 16#08#),
      2759 => to_slv(opcode_type, 16#0E#),
      2760 => to_slv(opcode_type, 16#0F#),
      2761 => to_slv(opcode_type, 16#C1#),
      2762 => to_slv(opcode_type, 16#0A#),
      2763 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#06#),
      2785 => to_slv(opcode_type, 16#02#),
      2786 => to_slv(opcode_type, 16#05#),
      2787 => to_slv(opcode_type, 16#06#),
      2788 => to_slv(opcode_type, 16#38#),
      2789 => to_slv(opcode_type, 16#5B#),
      2790 => to_slv(opcode_type, 16#05#),
      2791 => to_slv(opcode_type, 16#01#),
      2792 => to_slv(opcode_type, 16#08#),
      2793 => to_slv(opcode_type, 16#0A#),
      2794 => to_slv(opcode_type, 16#10#),
      2795 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#03#),
      2817 => to_slv(opcode_type, 16#08#),
      2818 => to_slv(opcode_type, 16#09#),
      2819 => to_slv(opcode_type, 16#08#),
      2820 => to_slv(opcode_type, 16#10#),
      2821 => to_slv(opcode_type, 16#0A#),
      2822 => to_slv(opcode_type, 16#05#),
      2823 => to_slv(opcode_type, 16#EA#),
      2824 => to_slv(opcode_type, 16#01#),
      2825 => to_slv(opcode_type, 16#03#),
      2826 => to_slv(opcode_type, 16#0E#),
      2827 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#03#),
      2849 => to_slv(opcode_type, 16#06#),
      2850 => to_slv(opcode_type, 16#07#),
      2851 => to_slv(opcode_type, 16#01#),
      2852 => to_slv(opcode_type, 16#0F#),
      2853 => to_slv(opcode_type, 16#06#),
      2854 => to_slv(opcode_type, 16#0F#),
      2855 => to_slv(opcode_type, 16#0C#),
      2856 => to_slv(opcode_type, 16#05#),
      2857 => to_slv(opcode_type, 16#02#),
      2858 => to_slv(opcode_type, 16#0F#),
      2859 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#04#),
      2881 => to_slv(opcode_type, 16#08#),
      2882 => to_slv(opcode_type, 16#01#),
      2883 => to_slv(opcode_type, 16#04#),
      2884 => to_slv(opcode_type, 16#79#),
      2885 => to_slv(opcode_type, 16#09#),
      2886 => to_slv(opcode_type, 16#01#),
      2887 => to_slv(opcode_type, 16#1C#),
      2888 => to_slv(opcode_type, 16#06#),
      2889 => to_slv(opcode_type, 16#0A#),
      2890 => to_slv(opcode_type, 16#11#),
      2891 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#04#),
      2913 => to_slv(opcode_type, 16#09#),
      2914 => to_slv(opcode_type, 16#03#),
      2915 => to_slv(opcode_type, 16#08#),
      2916 => to_slv(opcode_type, 16#11#),
      2917 => to_slv(opcode_type, 16#11#),
      2918 => to_slv(opcode_type, 16#09#),
      2919 => to_slv(opcode_type, 16#08#),
      2920 => to_slv(opcode_type, 16#0A#),
      2921 => to_slv(opcode_type, 16#10#),
      2922 => to_slv(opcode_type, 16#10#),
      2923 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#03#),
      2945 => to_slv(opcode_type, 16#09#),
      2946 => to_slv(opcode_type, 16#08#),
      2947 => to_slv(opcode_type, 16#08#),
      2948 => to_slv(opcode_type, 16#9F#),
      2949 => to_slv(opcode_type, 16#0F#),
      2950 => to_slv(opcode_type, 16#04#),
      2951 => to_slv(opcode_type, 16#0A#),
      2952 => to_slv(opcode_type, 16#06#),
      2953 => to_slv(opcode_type, 16#0A#),
      2954 => to_slv(opcode_type, 16#11#),
      2955 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#09#),
      2977 => to_slv(opcode_type, 16#08#),
      2978 => to_slv(opcode_type, 16#01#),
      2979 => to_slv(opcode_type, 16#07#),
      2980 => to_slv(opcode_type, 16#64#),
      2981 => to_slv(opcode_type, 16#10#),
      2982 => to_slv(opcode_type, 16#05#),
      2983 => to_slv(opcode_type, 16#06#),
      2984 => to_slv(opcode_type, 16#0C#),
      2985 => to_slv(opcode_type, 16#11#),
      2986 => to_slv(opcode_type, 16#11#),
      2987 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#09#),
      3009 => to_slv(opcode_type, 16#03#),
      3010 => to_slv(opcode_type, 16#02#),
      3011 => to_slv(opcode_type, 16#08#),
      3012 => to_slv(opcode_type, 16#0F#),
      3013 => to_slv(opcode_type, 16#10#),
      3014 => to_slv(opcode_type, 16#09#),
      3015 => to_slv(opcode_type, 16#02#),
      3016 => to_slv(opcode_type, 16#02#),
      3017 => to_slv(opcode_type, 16#0E#),
      3018 => to_slv(opcode_type, 16#0B#),
      3019 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#07#),
      3041 => to_slv(opcode_type, 16#01#),
      3042 => to_slv(opcode_type, 16#05#),
      3043 => to_slv(opcode_type, 16#05#),
      3044 => to_slv(opcode_type, 16#EF#),
      3045 => to_slv(opcode_type, 16#03#),
      3046 => to_slv(opcode_type, 16#07#),
      3047 => to_slv(opcode_type, 16#03#),
      3048 => to_slv(opcode_type, 16#0C#),
      3049 => to_slv(opcode_type, 16#03#),
      3050 => to_slv(opcode_type, 16#11#),
      3051 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#01#),
      3073 => to_slv(opcode_type, 16#06#),
      3074 => to_slv(opcode_type, 16#07#),
      3075 => to_slv(opcode_type, 16#07#),
      3076 => to_slv(opcode_type, 16#0B#),
      3077 => to_slv(opcode_type, 16#0F#),
      3078 => to_slv(opcode_type, 16#08#),
      3079 => to_slv(opcode_type, 16#0D#),
      3080 => to_slv(opcode_type, 16#0F#),
      3081 => to_slv(opcode_type, 16#03#),
      3082 => to_slv(opcode_type, 16#11#),
      3083 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#04#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#04#),
      3107 => to_slv(opcode_type, 16#03#),
      3108 => to_slv(opcode_type, 16#0E#),
      3109 => to_slv(opcode_type, 16#07#),
      3110 => to_slv(opcode_type, 16#04#),
      3111 => to_slv(opcode_type, 16#11#),
      3112 => to_slv(opcode_type, 16#07#),
      3113 => to_slv(opcode_type, 16#0C#),
      3114 => to_slv(opcode_type, 16#11#),
      3115 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#09#),
      3137 => to_slv(opcode_type, 16#08#),
      3138 => to_slv(opcode_type, 16#04#),
      3139 => to_slv(opcode_type, 16#09#),
      3140 => to_slv(opcode_type, 16#0D#),
      3141 => to_slv(opcode_type, 16#0D#),
      3142 => to_slv(opcode_type, 16#06#),
      3143 => to_slv(opcode_type, 16#01#),
      3144 => to_slv(opcode_type, 16#0C#),
      3145 => to_slv(opcode_type, 16#0B#),
      3146 => to_slv(opcode_type, 16#0E#),
      3147 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#03#),
      3169 => to_slv(opcode_type, 16#07#),
      3170 => to_slv(opcode_type, 16#06#),
      3171 => to_slv(opcode_type, 16#04#),
      3172 => to_slv(opcode_type, 16#11#),
      3173 => to_slv(opcode_type, 16#09#),
      3174 => to_slv(opcode_type, 16#0E#),
      3175 => to_slv(opcode_type, 16#0B#),
      3176 => to_slv(opcode_type, 16#02#),
      3177 => to_slv(opcode_type, 16#01#),
      3178 => to_slv(opcode_type, 16#0F#),
      3179 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#07#),
      3201 => to_slv(opcode_type, 16#08#),
      3202 => to_slv(opcode_type, 16#08#),
      3203 => to_slv(opcode_type, 16#02#),
      3204 => to_slv(opcode_type, 16#B3#),
      3205 => to_slv(opcode_type, 16#03#),
      3206 => to_slv(opcode_type, 16#11#),
      3207 => to_slv(opcode_type, 16#02#),
      3208 => to_slv(opcode_type, 16#03#),
      3209 => to_slv(opcode_type, 16#10#),
      3210 => to_slv(opcode_type, 16#0B#),
      3211 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#04#),
      3233 => to_slv(opcode_type, 16#09#),
      3234 => to_slv(opcode_type, 16#04#),
      3235 => to_slv(opcode_type, 16#05#),
      3236 => to_slv(opcode_type, 16#0D#),
      3237 => to_slv(opcode_type, 16#09#),
      3238 => to_slv(opcode_type, 16#04#),
      3239 => to_slv(opcode_type, 16#0F#),
      3240 => to_slv(opcode_type, 16#09#),
      3241 => to_slv(opcode_type, 16#0B#),
      3242 => to_slv(opcode_type, 16#0A#),
      3243 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#03#),
      3265 => to_slv(opcode_type, 16#06#),
      3266 => to_slv(opcode_type, 16#06#),
      3267 => to_slv(opcode_type, 16#07#),
      3268 => to_slv(opcode_type, 16#40#),
      3269 => to_slv(opcode_type, 16#11#),
      3270 => to_slv(opcode_type, 16#06#),
      3271 => to_slv(opcode_type, 16#0C#),
      3272 => to_slv(opcode_type, 16#0B#),
      3273 => to_slv(opcode_type, 16#01#),
      3274 => to_slv(opcode_type, 16#10#),
      3275 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#05#),
      3297 => to_slv(opcode_type, 16#07#),
      3298 => to_slv(opcode_type, 16#07#),
      3299 => to_slv(opcode_type, 16#09#),
      3300 => to_slv(opcode_type, 16#0B#),
      3301 => to_slv(opcode_type, 16#E6#),
      3302 => to_slv(opcode_type, 16#03#),
      3303 => to_slv(opcode_type, 16#0D#),
      3304 => to_slv(opcode_type, 16#01#),
      3305 => to_slv(opcode_type, 16#03#),
      3306 => to_slv(opcode_type, 16#FE#),
      3307 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#02#),
      3329 => to_slv(opcode_type, 16#07#),
      3330 => to_slv(opcode_type, 16#08#),
      3331 => to_slv(opcode_type, 16#01#),
      3332 => to_slv(opcode_type, 16#0F#),
      3333 => to_slv(opcode_type, 16#07#),
      3334 => to_slv(opcode_type, 16#0D#),
      3335 => to_slv(opcode_type, 16#0C#),
      3336 => to_slv(opcode_type, 16#03#),
      3337 => to_slv(opcode_type, 16#03#),
      3338 => to_slv(opcode_type, 16#60#),
      3339 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#05#),
      3361 => to_slv(opcode_type, 16#06#),
      3362 => to_slv(opcode_type, 16#04#),
      3363 => to_slv(opcode_type, 16#08#),
      3364 => to_slv(opcode_type, 16#B4#),
      3365 => to_slv(opcode_type, 16#0C#),
      3366 => to_slv(opcode_type, 16#08#),
      3367 => to_slv(opcode_type, 16#03#),
      3368 => to_slv(opcode_type, 16#0C#),
      3369 => to_slv(opcode_type, 16#01#),
      3370 => to_slv(opcode_type, 16#0C#),
      3371 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#06#),
      3393 => to_slv(opcode_type, 16#04#),
      3394 => to_slv(opcode_type, 16#04#),
      3395 => to_slv(opcode_type, 16#03#),
      3396 => to_slv(opcode_type, 16#0D#),
      3397 => to_slv(opcode_type, 16#03#),
      3398 => to_slv(opcode_type, 16#07#),
      3399 => to_slv(opcode_type, 16#03#),
      3400 => to_slv(opcode_type, 16#0F#),
      3401 => to_slv(opcode_type, 16#01#),
      3402 => to_slv(opcode_type, 16#0F#),
      3403 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#06#),
      3425 => to_slv(opcode_type, 16#08#),
      3426 => to_slv(opcode_type, 16#03#),
      3427 => to_slv(opcode_type, 16#08#),
      3428 => to_slv(opcode_type, 16#11#),
      3429 => to_slv(opcode_type, 16#10#),
      3430 => to_slv(opcode_type, 16#07#),
      3431 => to_slv(opcode_type, 16#01#),
      3432 => to_slv(opcode_type, 16#0C#),
      3433 => to_slv(opcode_type, 16#0C#),
      3434 => to_slv(opcode_type, 16#10#),
      3435 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#05#),
      3457 => to_slv(opcode_type, 16#08#),
      3458 => to_slv(opcode_type, 16#06#),
      3459 => to_slv(opcode_type, 16#06#),
      3460 => to_slv(opcode_type, 16#0D#),
      3461 => to_slv(opcode_type, 16#0B#),
      3462 => to_slv(opcode_type, 16#01#),
      3463 => to_slv(opcode_type, 16#B8#),
      3464 => to_slv(opcode_type, 16#05#),
      3465 => to_slv(opcode_type, 16#01#),
      3466 => to_slv(opcode_type, 16#0E#),
      3467 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#07#),
      3489 => to_slv(opcode_type, 16#05#),
      3490 => to_slv(opcode_type, 16#02#),
      3491 => to_slv(opcode_type, 16#02#),
      3492 => to_slv(opcode_type, 16#0D#),
      3493 => to_slv(opcode_type, 16#03#),
      3494 => to_slv(opcode_type, 16#08#),
      3495 => to_slv(opcode_type, 16#03#),
      3496 => to_slv(opcode_type, 16#0F#),
      3497 => to_slv(opcode_type, 16#03#),
      3498 => to_slv(opcode_type, 16#0D#),
      3499 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#08#),
      3521 => to_slv(opcode_type, 16#05#),
      3522 => to_slv(opcode_type, 16#03#),
      3523 => to_slv(opcode_type, 16#08#),
      3524 => to_slv(opcode_type, 16#0A#),
      3525 => to_slv(opcode_type, 16#0A#),
      3526 => to_slv(opcode_type, 16#07#),
      3527 => to_slv(opcode_type, 16#08#),
      3528 => to_slv(opcode_type, 16#0A#),
      3529 => to_slv(opcode_type, 16#0B#),
      3530 => to_slv(opcode_type, 16#0E#),
      3531 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#04#),
      3553 => to_slv(opcode_type, 16#07#),
      3554 => to_slv(opcode_type, 16#07#),
      3555 => to_slv(opcode_type, 16#06#),
      3556 => to_slv(opcode_type, 16#0C#),
      3557 => to_slv(opcode_type, 16#11#),
      3558 => to_slv(opcode_type, 16#06#),
      3559 => to_slv(opcode_type, 16#11#),
      3560 => to_slv(opcode_type, 16#0B#),
      3561 => to_slv(opcode_type, 16#02#),
      3562 => to_slv(opcode_type, 16#0F#),
      3563 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#01#),
      3585 => to_slv(opcode_type, 16#08#),
      3586 => to_slv(opcode_type, 16#08#),
      3587 => to_slv(opcode_type, 16#04#),
      3588 => to_slv(opcode_type, 16#0B#),
      3589 => to_slv(opcode_type, 16#09#),
      3590 => to_slv(opcode_type, 16#0C#),
      3591 => to_slv(opcode_type, 16#0C#),
      3592 => to_slv(opcode_type, 16#04#),
      3593 => to_slv(opcode_type, 16#02#),
      3594 => to_slv(opcode_type, 16#0C#),
      3595 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#09#),
      3617 => to_slv(opcode_type, 16#05#),
      3618 => to_slv(opcode_type, 16#01#),
      3619 => to_slv(opcode_type, 16#07#),
      3620 => to_slv(opcode_type, 16#0C#),
      3621 => to_slv(opcode_type, 16#70#),
      3622 => to_slv(opcode_type, 16#06#),
      3623 => to_slv(opcode_type, 16#07#),
      3624 => to_slv(opcode_type, 16#0E#),
      3625 => to_slv(opcode_type, 16#11#),
      3626 => to_slv(opcode_type, 16#0D#),
      3627 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#03#),
      3649 => to_slv(opcode_type, 16#08#),
      3650 => to_slv(opcode_type, 16#09#),
      3651 => to_slv(opcode_type, 16#02#),
      3652 => to_slv(opcode_type, 16#10#),
      3653 => to_slv(opcode_type, 16#07#),
      3654 => to_slv(opcode_type, 16#0C#),
      3655 => to_slv(opcode_type, 16#0B#),
      3656 => to_slv(opcode_type, 16#04#),
      3657 => to_slv(opcode_type, 16#04#),
      3658 => to_slv(opcode_type, 16#0A#),
      3659 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#06#),
      3681 => to_slv(opcode_type, 16#09#),
      3682 => to_slv(opcode_type, 16#01#),
      3683 => to_slv(opcode_type, 16#07#),
      3684 => to_slv(opcode_type, 16#11#),
      3685 => to_slv(opcode_type, 16#0A#),
      3686 => to_slv(opcode_type, 16#04#),
      3687 => to_slv(opcode_type, 16#06#),
      3688 => to_slv(opcode_type, 16#0B#),
      3689 => to_slv(opcode_type, 16#0F#),
      3690 => to_slv(opcode_type, 16#0A#),
      3691 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#01#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#04#),
      3715 => to_slv(opcode_type, 16#03#),
      3716 => to_slv(opcode_type, 16#0B#),
      3717 => to_slv(opcode_type, 16#08#),
      3718 => to_slv(opcode_type, 16#05#),
      3719 => to_slv(opcode_type, 16#11#),
      3720 => to_slv(opcode_type, 16#09#),
      3721 => to_slv(opcode_type, 16#0F#),
      3722 => to_slv(opcode_type, 16#0F#),
      3723 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#07#),
      3745 => to_slv(opcode_type, 16#01#),
      3746 => to_slv(opcode_type, 16#09#),
      3747 => to_slv(opcode_type, 16#09#),
      3748 => to_slv(opcode_type, 16#0F#),
      3749 => to_slv(opcode_type, 16#0C#),
      3750 => to_slv(opcode_type, 16#04#),
      3751 => to_slv(opcode_type, 16#0C#),
      3752 => to_slv(opcode_type, 16#08#),
      3753 => to_slv(opcode_type, 16#0E#),
      3754 => to_slv(opcode_type, 16#0D#),
      3755 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#02#),
      3777 => to_slv(opcode_type, 16#06#),
      3778 => to_slv(opcode_type, 16#04#),
      3779 => to_slv(opcode_type, 16#08#),
      3780 => to_slv(opcode_type, 16#11#),
      3781 => to_slv(opcode_type, 16#9D#),
      3782 => to_slv(opcode_type, 16#06#),
      3783 => to_slv(opcode_type, 16#08#),
      3784 => to_slv(opcode_type, 16#11#),
      3785 => to_slv(opcode_type, 16#0A#),
      3786 => to_slv(opcode_type, 16#0B#),
      3787 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#04#),
      3809 => to_slv(opcode_type, 16#09#),
      3810 => to_slv(opcode_type, 16#08#),
      3811 => to_slv(opcode_type, 16#04#),
      3812 => to_slv(opcode_type, 16#0C#),
      3813 => to_slv(opcode_type, 16#02#),
      3814 => to_slv(opcode_type, 16#0D#),
      3815 => to_slv(opcode_type, 16#03#),
      3816 => to_slv(opcode_type, 16#08#),
      3817 => to_slv(opcode_type, 16#0A#),
      3818 => to_slv(opcode_type, 16#F8#),
      3819 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#06#),
      3841 => to_slv(opcode_type, 16#08#),
      3842 => to_slv(opcode_type, 16#02#),
      3843 => to_slv(opcode_type, 16#02#),
      3844 => to_slv(opcode_type, 16#0F#),
      3845 => to_slv(opcode_type, 16#03#),
      3846 => to_slv(opcode_type, 16#07#),
      3847 => to_slv(opcode_type, 16#0E#),
      3848 => to_slv(opcode_type, 16#11#),
      3849 => to_slv(opcode_type, 16#04#),
      3850 => to_slv(opcode_type, 16#0C#),
      3851 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#06#),
      3873 => to_slv(opcode_type, 16#04#),
      3874 => to_slv(opcode_type, 16#04#),
      3875 => to_slv(opcode_type, 16#04#),
      3876 => to_slv(opcode_type, 16#0B#),
      3877 => to_slv(opcode_type, 16#05#),
      3878 => to_slv(opcode_type, 16#07#),
      3879 => to_slv(opcode_type, 16#04#),
      3880 => to_slv(opcode_type, 16#0C#),
      3881 => to_slv(opcode_type, 16#05#),
      3882 => to_slv(opcode_type, 16#0B#),
      3883 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#02#),
      3905 => to_slv(opcode_type, 16#07#),
      3906 => to_slv(opcode_type, 16#04#),
      3907 => to_slv(opcode_type, 16#08#),
      3908 => to_slv(opcode_type, 16#0C#),
      3909 => to_slv(opcode_type, 16#0A#),
      3910 => to_slv(opcode_type, 16#06#),
      3911 => to_slv(opcode_type, 16#06#),
      3912 => to_slv(opcode_type, 16#CE#),
      3913 => to_slv(opcode_type, 16#11#),
      3914 => to_slv(opcode_type, 16#0E#),
      3915 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#04#),
      3937 => to_slv(opcode_type, 16#09#),
      3938 => to_slv(opcode_type, 16#03#),
      3939 => to_slv(opcode_type, 16#02#),
      3940 => to_slv(opcode_type, 16#10#),
      3941 => to_slv(opcode_type, 16#07#),
      3942 => to_slv(opcode_type, 16#03#),
      3943 => to_slv(opcode_type, 16#10#),
      3944 => to_slv(opcode_type, 16#06#),
      3945 => to_slv(opcode_type, 16#0A#),
      3946 => to_slv(opcode_type, 16#0B#),
      3947 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#01#),
      3969 => to_slv(opcode_type, 16#07#),
      3970 => to_slv(opcode_type, 16#07#),
      3971 => to_slv(opcode_type, 16#08#),
      3972 => to_slv(opcode_type, 16#0A#),
      3973 => to_slv(opcode_type, 16#10#),
      3974 => to_slv(opcode_type, 16#04#),
      3975 => to_slv(opcode_type, 16#FA#),
      3976 => to_slv(opcode_type, 16#02#),
      3977 => to_slv(opcode_type, 16#02#),
      3978 => to_slv(opcode_type, 16#0A#),
      3979 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#04#),
      4001 => to_slv(opcode_type, 16#06#),
      4002 => to_slv(opcode_type, 16#06#),
      4003 => to_slv(opcode_type, 16#07#),
      4004 => to_slv(opcode_type, 16#0B#),
      4005 => to_slv(opcode_type, 16#10#),
      4006 => to_slv(opcode_type, 16#07#),
      4007 => to_slv(opcode_type, 16#11#),
      4008 => to_slv(opcode_type, 16#0B#),
      4009 => to_slv(opcode_type, 16#03#),
      4010 => to_slv(opcode_type, 16#0F#),
      4011 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#09#),
      4033 => to_slv(opcode_type, 16#07#),
      4034 => to_slv(opcode_type, 16#01#),
      4035 => to_slv(opcode_type, 16#02#),
      4036 => to_slv(opcode_type, 16#0A#),
      4037 => to_slv(opcode_type, 16#08#),
      4038 => to_slv(opcode_type, 16#09#),
      4039 => to_slv(opcode_type, 16#10#),
      4040 => to_slv(opcode_type, 16#10#),
      4041 => to_slv(opcode_type, 16#0E#),
      4042 => to_slv(opcode_type, 16#A7#),
      4043 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#04#),
      4066 => to_slv(opcode_type, 16#08#),
      4067 => to_slv(opcode_type, 16#03#),
      4068 => to_slv(opcode_type, 16#10#),
      4069 => to_slv(opcode_type, 16#03#),
      4070 => to_slv(opcode_type, 16#0D#),
      4071 => to_slv(opcode_type, 16#02#),
      4072 => to_slv(opcode_type, 16#06#),
      4073 => to_slv(opcode_type, 16#10#),
      4074 => to_slv(opcode_type, 16#0E#),
      4075 to 4095 => (others => '0')
  ),

    -- Bin `12`...
    11 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#09#),
      1 => to_slv(opcode_type, 16#04#),
      2 => to_slv(opcode_type, 16#01#),
      3 => to_slv(opcode_type, 16#03#),
      4 => to_slv(opcode_type, 16#0E#),
      5 => to_slv(opcode_type, 16#03#),
      6 => to_slv(opcode_type, 16#06#),
      7 => to_slv(opcode_type, 16#04#),
      8 => to_slv(opcode_type, 16#11#),
      9 => to_slv(opcode_type, 16#07#),
      10 => to_slv(opcode_type, 16#0D#),
      11 => to_slv(opcode_type, 16#0F#),
      12 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#04#),
      33 => to_slv(opcode_type, 16#09#),
      34 => to_slv(opcode_type, 16#02#),
      35 => to_slv(opcode_type, 16#01#),
      36 => to_slv(opcode_type, 16#0F#),
      37 => to_slv(opcode_type, 16#07#),
      38 => to_slv(opcode_type, 16#07#),
      39 => to_slv(opcode_type, 16#56#),
      40 => to_slv(opcode_type, 16#10#),
      41 => to_slv(opcode_type, 16#06#),
      42 => to_slv(opcode_type, 16#0B#),
      43 => to_slv(opcode_type, 16#11#),
      44 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#05#),
      65 => to_slv(opcode_type, 16#06#),
      66 => to_slv(opcode_type, 16#03#),
      67 => to_slv(opcode_type, 16#01#),
      68 => to_slv(opcode_type, 16#0A#),
      69 => to_slv(opcode_type, 16#06#),
      70 => to_slv(opcode_type, 16#06#),
      71 => to_slv(opcode_type, 16#11#),
      72 => to_slv(opcode_type, 16#0A#),
      73 => to_slv(opcode_type, 16#07#),
      74 => to_slv(opcode_type, 16#0B#),
      75 => to_slv(opcode_type, 16#0C#),
      76 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#07#),
      97 => to_slv(opcode_type, 16#03#),
      98 => to_slv(opcode_type, 16#07#),
      99 => to_slv(opcode_type, 16#03#),
      100 => to_slv(opcode_type, 16#0E#),
      101 => to_slv(opcode_type, 16#09#),
      102 => to_slv(opcode_type, 16#0A#),
      103 => to_slv(opcode_type, 16#10#),
      104 => to_slv(opcode_type, 16#05#),
      105 => to_slv(opcode_type, 16#06#),
      106 => to_slv(opcode_type, 16#0A#),
      107 => to_slv(opcode_type, 16#0F#),
      108 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#01#),
      129 => to_slv(opcode_type, 16#08#),
      130 => to_slv(opcode_type, 16#04#),
      131 => to_slv(opcode_type, 16#04#),
      132 => to_slv(opcode_type, 16#0B#),
      133 => to_slv(opcode_type, 16#07#),
      134 => to_slv(opcode_type, 16#07#),
      135 => to_slv(opcode_type, 16#10#),
      136 => to_slv(opcode_type, 16#B2#),
      137 => to_slv(opcode_type, 16#09#),
      138 => to_slv(opcode_type, 16#4B#),
      139 => to_slv(opcode_type, 16#0B#),
      140 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#05#),
      161 => to_slv(opcode_type, 16#08#),
      162 => to_slv(opcode_type, 16#06#),
      163 => to_slv(opcode_type, 16#05#),
      164 => to_slv(opcode_type, 16#0C#),
      165 => to_slv(opcode_type, 16#09#),
      166 => to_slv(opcode_type, 16#0F#),
      167 => to_slv(opcode_type, 16#0A#),
      168 => to_slv(opcode_type, 16#05#),
      169 => to_slv(opcode_type, 16#07#),
      170 => to_slv(opcode_type, 16#0D#),
      171 => to_slv(opcode_type, 16#0F#),
      172 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#08#),
      193 => to_slv(opcode_type, 16#08#),
      194 => to_slv(opcode_type, 16#05#),
      195 => to_slv(opcode_type, 16#02#),
      196 => to_slv(opcode_type, 16#0B#),
      197 => to_slv(opcode_type, 16#01#),
      198 => to_slv(opcode_type, 16#07#),
      199 => to_slv(opcode_type, 16#10#),
      200 => to_slv(opcode_type, 16#0B#),
      201 => to_slv(opcode_type, 16#03#),
      202 => to_slv(opcode_type, 16#04#),
      203 => to_slv(opcode_type, 16#0E#),
      204 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#08#),
      225 => to_slv(opcode_type, 16#03#),
      226 => to_slv(opcode_type, 16#02#),
      227 => to_slv(opcode_type, 16#05#),
      228 => to_slv(opcode_type, 16#0F#),
      229 => to_slv(opcode_type, 16#06#),
      230 => to_slv(opcode_type, 16#02#),
      231 => to_slv(opcode_type, 16#03#),
      232 => to_slv(opcode_type, 16#0F#),
      233 => to_slv(opcode_type, 16#04#),
      234 => to_slv(opcode_type, 16#05#),
      235 => to_slv(opcode_type, 16#10#),
      236 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#04#),
      257 => to_slv(opcode_type, 16#07#),
      258 => to_slv(opcode_type, 16#01#),
      259 => to_slv(opcode_type, 16#05#),
      260 => to_slv(opcode_type, 16#0A#),
      261 => to_slv(opcode_type, 16#08#),
      262 => to_slv(opcode_type, 16#08#),
      263 => to_slv(opcode_type, 16#0C#),
      264 => to_slv(opcode_type, 16#5D#),
      265 => to_slv(opcode_type, 16#07#),
      266 => to_slv(opcode_type, 16#18#),
      267 => to_slv(opcode_type, 16#11#),
      268 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#01#),
      289 => to_slv(opcode_type, 16#06#),
      290 => to_slv(opcode_type, 16#07#),
      291 => to_slv(opcode_type, 16#01#),
      292 => to_slv(opcode_type, 16#0A#),
      293 => to_slv(opcode_type, 16#04#),
      294 => to_slv(opcode_type, 16#0B#),
      295 => to_slv(opcode_type, 16#07#),
      296 => to_slv(opcode_type, 16#07#),
      297 => to_slv(opcode_type, 16#6E#),
      298 => to_slv(opcode_type, 16#11#),
      299 => to_slv(opcode_type, 16#0D#),
      300 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#09#),
      321 => to_slv(opcode_type, 16#06#),
      322 => to_slv(opcode_type, 16#08#),
      323 => to_slv(opcode_type, 16#02#),
      324 => to_slv(opcode_type, 16#0A#),
      325 => to_slv(opcode_type, 16#04#),
      326 => to_slv(opcode_type, 16#0F#),
      327 => to_slv(opcode_type, 16#01#),
      328 => to_slv(opcode_type, 16#04#),
      329 => to_slv(opcode_type, 16#0B#),
      330 => to_slv(opcode_type, 16#05#),
      331 => to_slv(opcode_type, 16#19#),
      332 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#09#),
      353 => to_slv(opcode_type, 16#08#),
      354 => to_slv(opcode_type, 16#05#),
      355 => to_slv(opcode_type, 16#09#),
      356 => to_slv(opcode_type, 16#10#),
      357 => to_slv(opcode_type, 16#0D#),
      358 => to_slv(opcode_type, 16#05#),
      359 => to_slv(opcode_type, 16#09#),
      360 => to_slv(opcode_type, 16#10#),
      361 => to_slv(opcode_type, 16#11#),
      362 => to_slv(opcode_type, 16#03#),
      363 => to_slv(opcode_type, 16#0B#),
      364 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#04#),
      385 => to_slv(opcode_type, 16#08#),
      386 => to_slv(opcode_type, 16#02#),
      387 => to_slv(opcode_type, 16#04#),
      388 => to_slv(opcode_type, 16#0B#),
      389 => to_slv(opcode_type, 16#08#),
      390 => to_slv(opcode_type, 16#09#),
      391 => to_slv(opcode_type, 16#11#),
      392 => to_slv(opcode_type, 16#0F#),
      393 => to_slv(opcode_type, 16#08#),
      394 => to_slv(opcode_type, 16#0E#),
      395 => to_slv(opcode_type, 16#0B#),
      396 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#08#),
      417 => to_slv(opcode_type, 16#08#),
      418 => to_slv(opcode_type, 16#05#),
      419 => to_slv(opcode_type, 16#08#),
      420 => to_slv(opcode_type, 16#10#),
      421 => to_slv(opcode_type, 16#10#),
      422 => to_slv(opcode_type, 16#03#),
      423 => to_slv(opcode_type, 16#02#),
      424 => to_slv(opcode_type, 16#0F#),
      425 => to_slv(opcode_type, 16#07#),
      426 => to_slv(opcode_type, 16#0D#),
      427 => to_slv(opcode_type, 16#0F#),
      428 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#09#),
      449 => to_slv(opcode_type, 16#06#),
      450 => to_slv(opcode_type, 16#09#),
      451 => to_slv(opcode_type, 16#07#),
      452 => to_slv(opcode_type, 16#11#),
      453 => to_slv(opcode_type, 16#0B#),
      454 => to_slv(opcode_type, 16#03#),
      455 => to_slv(opcode_type, 16#0D#),
      456 => to_slv(opcode_type, 16#06#),
      457 => to_slv(opcode_type, 16#0D#),
      458 => to_slv(opcode_type, 16#0C#),
      459 => to_slv(opcode_type, 16#0F#),
      460 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#05#),
      481 => to_slv(opcode_type, 16#07#),
      482 => to_slv(opcode_type, 16#02#),
      483 => to_slv(opcode_type, 16#02#),
      484 => to_slv(opcode_type, 16#0F#),
      485 => to_slv(opcode_type, 16#07#),
      486 => to_slv(opcode_type, 16#08#),
      487 => to_slv(opcode_type, 16#0A#),
      488 => to_slv(opcode_type, 16#0E#),
      489 => to_slv(opcode_type, 16#06#),
      490 => to_slv(opcode_type, 16#0B#),
      491 => to_slv(opcode_type, 16#10#),
      492 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#08#),
      513 => to_slv(opcode_type, 16#01#),
      514 => to_slv(opcode_type, 16#01#),
      515 => to_slv(opcode_type, 16#09#),
      516 => to_slv(opcode_type, 16#D4#),
      517 => to_slv(opcode_type, 16#0A#),
      518 => to_slv(opcode_type, 16#03#),
      519 => to_slv(opcode_type, 16#09#),
      520 => to_slv(opcode_type, 16#06#),
      521 => to_slv(opcode_type, 16#0C#),
      522 => to_slv(opcode_type, 16#0A#),
      523 => to_slv(opcode_type, 16#0B#),
      524 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#08#),
      545 => to_slv(opcode_type, 16#01#),
      546 => to_slv(opcode_type, 16#04#),
      547 => to_slv(opcode_type, 16#06#),
      548 => to_slv(opcode_type, 16#DC#),
      549 => to_slv(opcode_type, 16#0D#),
      550 => to_slv(opcode_type, 16#09#),
      551 => to_slv(opcode_type, 16#07#),
      552 => to_slv(opcode_type, 16#05#),
      553 => to_slv(opcode_type, 16#0A#),
      554 => to_slv(opcode_type, 16#0A#),
      555 => to_slv(opcode_type, 16#0D#),
      556 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#01#),
      577 => to_slv(opcode_type, 16#09#),
      578 => to_slv(opcode_type, 16#05#),
      579 => to_slv(opcode_type, 16#09#),
      580 => to_slv(opcode_type, 16#0E#),
      581 => to_slv(opcode_type, 16#0F#),
      582 => to_slv(opcode_type, 16#08#),
      583 => to_slv(opcode_type, 16#04#),
      584 => to_slv(opcode_type, 16#0E#),
      585 => to_slv(opcode_type, 16#09#),
      586 => to_slv(opcode_type, 16#0B#),
      587 => to_slv(opcode_type, 16#0E#),
      588 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#08#),
      609 => to_slv(opcode_type, 16#02#),
      610 => to_slv(opcode_type, 16#01#),
      611 => to_slv(opcode_type, 16#08#),
      612 => to_slv(opcode_type, 16#10#),
      613 => to_slv(opcode_type, 16#0E#),
      614 => to_slv(opcode_type, 16#08#),
      615 => to_slv(opcode_type, 16#06#),
      616 => to_slv(opcode_type, 16#05#),
      617 => to_slv(opcode_type, 16#BD#),
      618 => to_slv(opcode_type, 16#5F#),
      619 => to_slv(opcode_type, 16#0E#),
      620 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#05#),
      641 => to_slv(opcode_type, 16#09#),
      642 => to_slv(opcode_type, 16#07#),
      643 => to_slv(opcode_type, 16#05#),
      644 => to_slv(opcode_type, 16#10#),
      645 => to_slv(opcode_type, 16#07#),
      646 => to_slv(opcode_type, 16#11#),
      647 => to_slv(opcode_type, 16#0A#),
      648 => to_slv(opcode_type, 16#08#),
      649 => to_slv(opcode_type, 16#05#),
      650 => to_slv(opcode_type, 16#10#),
      651 => to_slv(opcode_type, 16#11#),
      652 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#05#),
      673 => to_slv(opcode_type, 16#06#),
      674 => to_slv(opcode_type, 16#06#),
      675 => to_slv(opcode_type, 16#09#),
      676 => to_slv(opcode_type, 16#11#),
      677 => to_slv(opcode_type, 16#0D#),
      678 => to_slv(opcode_type, 16#05#),
      679 => to_slv(opcode_type, 16#0D#),
      680 => to_slv(opcode_type, 16#01#),
      681 => to_slv(opcode_type, 16#06#),
      682 => to_slv(opcode_type, 16#0B#),
      683 => to_slv(opcode_type, 16#10#),
      684 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#06#),
      705 => to_slv(opcode_type, 16#08#),
      706 => to_slv(opcode_type, 16#02#),
      707 => to_slv(opcode_type, 16#05#),
      708 => to_slv(opcode_type, 16#0A#),
      709 => to_slv(opcode_type, 16#09#),
      710 => to_slv(opcode_type, 16#05#),
      711 => to_slv(opcode_type, 16#0C#),
      712 => to_slv(opcode_type, 16#02#),
      713 => to_slv(opcode_type, 16#10#),
      714 => to_slv(opcode_type, 16#03#),
      715 => to_slv(opcode_type, 16#0A#),
      716 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#04#),
      737 => to_slv(opcode_type, 16#07#),
      738 => to_slv(opcode_type, 16#08#),
      739 => to_slv(opcode_type, 16#07#),
      740 => to_slv(opcode_type, 16#0C#),
      741 => to_slv(opcode_type, 16#0C#),
      742 => to_slv(opcode_type, 16#03#),
      743 => to_slv(opcode_type, 16#11#),
      744 => to_slv(opcode_type, 16#08#),
      745 => to_slv(opcode_type, 16#05#),
      746 => to_slv(opcode_type, 16#10#),
      747 => to_slv(opcode_type, 16#11#),
      748 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#06#),
      769 => to_slv(opcode_type, 16#03#),
      770 => to_slv(opcode_type, 16#05#),
      771 => to_slv(opcode_type, 16#03#),
      772 => to_slv(opcode_type, 16#11#),
      773 => to_slv(opcode_type, 16#05#),
      774 => to_slv(opcode_type, 16#09#),
      775 => to_slv(opcode_type, 16#01#),
      776 => to_slv(opcode_type, 16#0F#),
      777 => to_slv(opcode_type, 16#06#),
      778 => to_slv(opcode_type, 16#0B#),
      779 => to_slv(opcode_type, 16#10#),
      780 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#03#),
      801 => to_slv(opcode_type, 16#09#),
      802 => to_slv(opcode_type, 16#02#),
      803 => to_slv(opcode_type, 16#05#),
      804 => to_slv(opcode_type, 16#0C#),
      805 => to_slv(opcode_type, 16#08#),
      806 => to_slv(opcode_type, 16#06#),
      807 => to_slv(opcode_type, 16#0E#),
      808 => to_slv(opcode_type, 16#0C#),
      809 => to_slv(opcode_type, 16#09#),
      810 => to_slv(opcode_type, 16#8B#),
      811 => to_slv(opcode_type, 16#0F#),
      812 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#05#),
      833 => to_slv(opcode_type, 16#07#),
      834 => to_slv(opcode_type, 16#08#),
      835 => to_slv(opcode_type, 16#03#),
      836 => to_slv(opcode_type, 16#10#),
      837 => to_slv(opcode_type, 16#02#),
      838 => to_slv(opcode_type, 16#0F#),
      839 => to_slv(opcode_type, 16#08#),
      840 => to_slv(opcode_type, 16#05#),
      841 => to_slv(opcode_type, 16#0E#),
      842 => to_slv(opcode_type, 16#01#),
      843 => to_slv(opcode_type, 16#0A#),
      844 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#01#),
      865 => to_slv(opcode_type, 16#09#),
      866 => to_slv(opcode_type, 16#02#),
      867 => to_slv(opcode_type, 16#01#),
      868 => to_slv(opcode_type, 16#CD#),
      869 => to_slv(opcode_type, 16#07#),
      870 => to_slv(opcode_type, 16#07#),
      871 => to_slv(opcode_type, 16#0E#),
      872 => to_slv(opcode_type, 16#11#),
      873 => to_slv(opcode_type, 16#06#),
      874 => to_slv(opcode_type, 16#0E#),
      875 => to_slv(opcode_type, 16#11#),
      876 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#07#),
      898 => to_slv(opcode_type, 16#02#),
      899 => to_slv(opcode_type, 16#01#),
      900 => to_slv(opcode_type, 16#11#),
      901 => to_slv(opcode_type, 16#07#),
      902 => to_slv(opcode_type, 16#09#),
      903 => to_slv(opcode_type, 16#76#),
      904 => to_slv(opcode_type, 16#11#),
      905 => to_slv(opcode_type, 16#03#),
      906 => to_slv(opcode_type, 16#0A#),
      907 => to_slv(opcode_type, 16#0F#),
      908 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#04#),
      929 => to_slv(opcode_type, 16#07#),
      930 => to_slv(opcode_type, 16#06#),
      931 => to_slv(opcode_type, 16#07#),
      932 => to_slv(opcode_type, 16#11#),
      933 => to_slv(opcode_type, 16#0F#),
      934 => to_slv(opcode_type, 16#05#),
      935 => to_slv(opcode_type, 16#0E#),
      936 => to_slv(opcode_type, 16#06#),
      937 => to_slv(opcode_type, 16#05#),
      938 => to_slv(opcode_type, 16#3F#),
      939 => to_slv(opcode_type, 16#0D#),
      940 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#01#),
      961 => to_slv(opcode_type, 16#08#),
      962 => to_slv(opcode_type, 16#09#),
      963 => to_slv(opcode_type, 16#05#),
      964 => to_slv(opcode_type, 16#1C#),
      965 => to_slv(opcode_type, 16#02#),
      966 => to_slv(opcode_type, 16#73#),
      967 => to_slv(opcode_type, 16#06#),
      968 => to_slv(opcode_type, 16#01#),
      969 => to_slv(opcode_type, 16#0F#),
      970 => to_slv(opcode_type, 16#02#),
      971 => to_slv(opcode_type, 16#0F#),
      972 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#05#),
      993 => to_slv(opcode_type, 16#06#),
      994 => to_slv(opcode_type, 16#09#),
      995 => to_slv(opcode_type, 16#03#),
      996 => to_slv(opcode_type, 16#0B#),
      997 => to_slv(opcode_type, 16#02#),
      998 => to_slv(opcode_type, 16#0D#),
      999 => to_slv(opcode_type, 16#09#),
      1000 => to_slv(opcode_type, 16#09#),
      1001 => to_slv(opcode_type, 16#C5#),
      1002 => to_slv(opcode_type, 16#0F#),
      1003 => to_slv(opcode_type, 16#0F#),
      1004 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#07#),
      1025 => to_slv(opcode_type, 16#01#),
      1026 => to_slv(opcode_type, 16#03#),
      1027 => to_slv(opcode_type, 16#05#),
      1028 => to_slv(opcode_type, 16#0C#),
      1029 => to_slv(opcode_type, 16#01#),
      1030 => to_slv(opcode_type, 16#06#),
      1031 => to_slv(opcode_type, 16#06#),
      1032 => to_slv(opcode_type, 16#0C#),
      1033 => to_slv(opcode_type, 16#0A#),
      1034 => to_slv(opcode_type, 16#01#),
      1035 => to_slv(opcode_type, 16#0F#),
      1036 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#04#),
      1057 => to_slv(opcode_type, 16#08#),
      1058 => to_slv(opcode_type, 16#02#),
      1059 => to_slv(opcode_type, 16#06#),
      1060 => to_slv(opcode_type, 16#46#),
      1061 => to_slv(opcode_type, 16#10#),
      1062 => to_slv(opcode_type, 16#07#),
      1063 => to_slv(opcode_type, 16#06#),
      1064 => to_slv(opcode_type, 16#0A#),
      1065 => to_slv(opcode_type, 16#0A#),
      1066 => to_slv(opcode_type, 16#01#),
      1067 => to_slv(opcode_type, 16#0B#),
      1068 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#09#),
      1089 => to_slv(opcode_type, 16#01#),
      1090 => to_slv(opcode_type, 16#06#),
      1091 => to_slv(opcode_type, 16#08#),
      1092 => to_slv(opcode_type, 16#0D#),
      1093 => to_slv(opcode_type, 16#10#),
      1094 => to_slv(opcode_type, 16#06#),
      1095 => to_slv(opcode_type, 16#0A#),
      1096 => to_slv(opcode_type, 16#11#),
      1097 => to_slv(opcode_type, 16#07#),
      1098 => to_slv(opcode_type, 16#0E#),
      1099 => to_slv(opcode_type, 16#C5#),
      1100 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#02#),
      1121 => to_slv(opcode_type, 16#06#),
      1122 => to_slv(opcode_type, 16#04#),
      1123 => to_slv(opcode_type, 16#04#),
      1124 => to_slv(opcode_type, 16#10#),
      1125 => to_slv(opcode_type, 16#06#),
      1126 => to_slv(opcode_type, 16#08#),
      1127 => to_slv(opcode_type, 16#11#),
      1128 => to_slv(opcode_type, 16#0C#),
      1129 => to_slv(opcode_type, 16#07#),
      1130 => to_slv(opcode_type, 16#11#),
      1131 => to_slv(opcode_type, 16#0D#),
      1132 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#07#),
      1153 => to_slv(opcode_type, 16#04#),
      1154 => to_slv(opcode_type, 16#09#),
      1155 => to_slv(opcode_type, 16#03#),
      1156 => to_slv(opcode_type, 16#0B#),
      1157 => to_slv(opcode_type, 16#08#),
      1158 => to_slv(opcode_type, 16#0A#),
      1159 => to_slv(opcode_type, 16#0B#),
      1160 => to_slv(opcode_type, 16#04#),
      1161 => to_slv(opcode_type, 16#01#),
      1162 => to_slv(opcode_type, 16#05#),
      1163 => to_slv(opcode_type, 16#0F#),
      1164 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#01#),
      1185 => to_slv(opcode_type, 16#09#),
      1186 => to_slv(opcode_type, 16#03#),
      1187 => to_slv(opcode_type, 16#07#),
      1188 => to_slv(opcode_type, 16#57#),
      1189 => to_slv(opcode_type, 16#0F#),
      1190 => to_slv(opcode_type, 16#06#),
      1191 => to_slv(opcode_type, 16#06#),
      1192 => to_slv(opcode_type, 16#4D#),
      1193 => to_slv(opcode_type, 16#0B#),
      1194 => to_slv(opcode_type, 16#01#),
      1195 => to_slv(opcode_type, 16#0E#),
      1196 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#02#),
      1217 => to_slv(opcode_type, 16#07#),
      1218 => to_slv(opcode_type, 16#06#),
      1219 => to_slv(opcode_type, 16#02#),
      1220 => to_slv(opcode_type, 16#0A#),
      1221 => to_slv(opcode_type, 16#07#),
      1222 => to_slv(opcode_type, 16#10#),
      1223 => to_slv(opcode_type, 16#0A#),
      1224 => to_slv(opcode_type, 16#04#),
      1225 => to_slv(opcode_type, 16#09#),
      1226 => to_slv(opcode_type, 16#0E#),
      1227 => to_slv(opcode_type, 16#0B#),
      1228 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#08#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#06#),
      1251 => to_slv(opcode_type, 16#06#),
      1252 => to_slv(opcode_type, 16#10#),
      1253 => to_slv(opcode_type, 16#0A#),
      1254 => to_slv(opcode_type, 16#03#),
      1255 => to_slv(opcode_type, 16#93#),
      1256 => to_slv(opcode_type, 16#07#),
      1257 => to_slv(opcode_type, 16#10#),
      1258 => to_slv(opcode_type, 16#0A#),
      1259 => to_slv(opcode_type, 16#0A#),
      1260 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#03#),
      1281 => to_slv(opcode_type, 16#08#),
      1282 => to_slv(opcode_type, 16#01#),
      1283 => to_slv(opcode_type, 16#06#),
      1284 => to_slv(opcode_type, 16#59#),
      1285 => to_slv(opcode_type, 16#11#),
      1286 => to_slv(opcode_type, 16#07#),
      1287 => to_slv(opcode_type, 16#03#),
      1288 => to_slv(opcode_type, 16#0A#),
      1289 => to_slv(opcode_type, 16#07#),
      1290 => to_slv(opcode_type, 16#0C#),
      1291 => to_slv(opcode_type, 16#0E#),
      1292 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#02#),
      1313 => to_slv(opcode_type, 16#06#),
      1314 => to_slv(opcode_type, 16#01#),
      1315 => to_slv(opcode_type, 16#07#),
      1316 => to_slv(opcode_type, 16#11#),
      1317 => to_slv(opcode_type, 16#0F#),
      1318 => to_slv(opcode_type, 16#07#),
      1319 => to_slv(opcode_type, 16#05#),
      1320 => to_slv(opcode_type, 16#D1#),
      1321 => to_slv(opcode_type, 16#09#),
      1322 => to_slv(opcode_type, 16#0A#),
      1323 => to_slv(opcode_type, 16#10#),
      1324 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#08#),
      1345 => to_slv(opcode_type, 16#07#),
      1346 => to_slv(opcode_type, 16#03#),
      1347 => to_slv(opcode_type, 16#05#),
      1348 => to_slv(opcode_type, 16#8D#),
      1349 => to_slv(opcode_type, 16#08#),
      1350 => to_slv(opcode_type, 16#02#),
      1351 => to_slv(opcode_type, 16#10#),
      1352 => to_slv(opcode_type, 16#05#),
      1353 => to_slv(opcode_type, 16#AE#),
      1354 => to_slv(opcode_type, 16#05#),
      1355 => to_slv(opcode_type, 16#0A#),
      1356 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#02#),
      1377 => to_slv(opcode_type, 16#07#),
      1378 => to_slv(opcode_type, 16#08#),
      1379 => to_slv(opcode_type, 16#05#),
      1380 => to_slv(opcode_type, 16#0E#),
      1381 => to_slv(opcode_type, 16#06#),
      1382 => to_slv(opcode_type, 16#0F#),
      1383 => to_slv(opcode_type, 16#59#),
      1384 => to_slv(opcode_type, 16#08#),
      1385 => to_slv(opcode_type, 16#01#),
      1386 => to_slv(opcode_type, 16#0F#),
      1387 => to_slv(opcode_type, 16#11#),
      1388 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#07#),
      1409 => to_slv(opcode_type, 16#08#),
      1410 => to_slv(opcode_type, 16#09#),
      1411 => to_slv(opcode_type, 16#02#),
      1412 => to_slv(opcode_type, 16#0F#),
      1413 => to_slv(opcode_type, 16#04#),
      1414 => to_slv(opcode_type, 16#0F#),
      1415 => to_slv(opcode_type, 16#08#),
      1416 => to_slv(opcode_type, 16#05#),
      1417 => to_slv(opcode_type, 16#CD#),
      1418 => to_slv(opcode_type, 16#64#),
      1419 => to_slv(opcode_type, 16#0A#),
      1420 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#02#),
      1441 => to_slv(opcode_type, 16#09#),
      1442 => to_slv(opcode_type, 16#09#),
      1443 => to_slv(opcode_type, 16#06#),
      1444 => to_slv(opcode_type, 16#11#),
      1445 => to_slv(opcode_type, 16#0A#),
      1446 => to_slv(opcode_type, 16#07#),
      1447 => to_slv(opcode_type, 16#0A#),
      1448 => to_slv(opcode_type, 16#10#),
      1449 => to_slv(opcode_type, 16#09#),
      1450 => to_slv(opcode_type, 16#0E#),
      1451 => to_slv(opcode_type, 16#0A#),
      1452 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#04#),
      1473 => to_slv(opcode_type, 16#06#),
      1474 => to_slv(opcode_type, 16#01#),
      1475 => to_slv(opcode_type, 16#08#),
      1476 => to_slv(opcode_type, 16#0B#),
      1477 => to_slv(opcode_type, 16#11#),
      1478 => to_slv(opcode_type, 16#06#),
      1479 => to_slv(opcode_type, 16#07#),
      1480 => to_slv(opcode_type, 16#11#),
      1481 => to_slv(opcode_type, 16#0B#),
      1482 => to_slv(opcode_type, 16#05#),
      1483 => to_slv(opcode_type, 16#0E#),
      1484 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#08#),
      1505 => to_slv(opcode_type, 16#06#),
      1506 => to_slv(opcode_type, 16#08#),
      1507 => to_slv(opcode_type, 16#09#),
      1508 => to_slv(opcode_type, 16#0F#),
      1509 => to_slv(opcode_type, 16#0C#),
      1510 => to_slv(opcode_type, 16#04#),
      1511 => to_slv(opcode_type, 16#0D#),
      1512 => to_slv(opcode_type, 16#08#),
      1513 => to_slv(opcode_type, 16#0C#),
      1514 => to_slv(opcode_type, 16#0E#),
      1515 => to_slv(opcode_type, 16#0A#),
      1516 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#05#),
      1537 => to_slv(opcode_type, 16#08#),
      1538 => to_slv(opcode_type, 16#02#),
      1539 => to_slv(opcode_type, 16#05#),
      1540 => to_slv(opcode_type, 16#0A#),
      1541 => to_slv(opcode_type, 16#08#),
      1542 => to_slv(opcode_type, 16#08#),
      1543 => to_slv(opcode_type, 16#0E#),
      1544 => to_slv(opcode_type, 16#0B#),
      1545 => to_slv(opcode_type, 16#07#),
      1546 => to_slv(opcode_type, 16#0E#),
      1547 => to_slv(opcode_type, 16#34#),
      1548 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#04#),
      1569 => to_slv(opcode_type, 16#06#),
      1570 => to_slv(opcode_type, 16#01#),
      1571 => to_slv(opcode_type, 16#07#),
      1572 => to_slv(opcode_type, 16#0D#),
      1573 => to_slv(opcode_type, 16#0E#),
      1574 => to_slv(opcode_type, 16#07#),
      1575 => to_slv(opcode_type, 16#01#),
      1576 => to_slv(opcode_type, 16#0A#),
      1577 => to_slv(opcode_type, 16#07#),
      1578 => to_slv(opcode_type, 16#CC#),
      1579 => to_slv(opcode_type, 16#0E#),
      1580 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#05#),
      1601 => to_slv(opcode_type, 16#09#),
      1602 => to_slv(opcode_type, 16#05#),
      1603 => to_slv(opcode_type, 16#01#),
      1604 => to_slv(opcode_type, 16#11#),
      1605 => to_slv(opcode_type, 16#09#),
      1606 => to_slv(opcode_type, 16#09#),
      1607 => to_slv(opcode_type, 16#0E#),
      1608 => to_slv(opcode_type, 16#0E#),
      1609 => to_slv(opcode_type, 16#06#),
      1610 => to_slv(opcode_type, 16#0B#),
      1611 => to_slv(opcode_type, 16#0E#),
      1612 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#04#),
      1633 => to_slv(opcode_type, 16#08#),
      1634 => to_slv(opcode_type, 16#09#),
      1635 => to_slv(opcode_type, 16#03#),
      1636 => to_slv(opcode_type, 16#10#),
      1637 => to_slv(opcode_type, 16#06#),
      1638 => to_slv(opcode_type, 16#10#),
      1639 => to_slv(opcode_type, 16#0A#),
      1640 => to_slv(opcode_type, 16#03#),
      1641 => to_slv(opcode_type, 16#06#),
      1642 => to_slv(opcode_type, 16#0B#),
      1643 => to_slv(opcode_type, 16#5A#),
      1644 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#04#),
      1666 => to_slv(opcode_type, 16#09#),
      1667 => to_slv(opcode_type, 16#07#),
      1668 => to_slv(opcode_type, 16#0E#),
      1669 => to_slv(opcode_type, 16#0C#),
      1670 => to_slv(opcode_type, 16#05#),
      1671 => to_slv(opcode_type, 16#11#),
      1672 => to_slv(opcode_type, 16#06#),
      1673 => to_slv(opcode_type, 16#04#),
      1674 => to_slv(opcode_type, 16#0D#),
      1675 => to_slv(opcode_type, 16#0B#),
      1676 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#02#),
      1697 => to_slv(opcode_type, 16#06#),
      1698 => to_slv(opcode_type, 16#01#),
      1699 => to_slv(opcode_type, 16#07#),
      1700 => to_slv(opcode_type, 16#0C#),
      1701 => to_slv(opcode_type, 16#10#),
      1702 => to_slv(opcode_type, 16#09#),
      1703 => to_slv(opcode_type, 16#07#),
      1704 => to_slv(opcode_type, 16#0C#),
      1705 => to_slv(opcode_type, 16#53#),
      1706 => to_slv(opcode_type, 16#05#),
      1707 => to_slv(opcode_type, 16#3A#),
      1708 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#09#),
      1729 => to_slv(opcode_type, 16#02#),
      1730 => to_slv(opcode_type, 16#07#),
      1731 => to_slv(opcode_type, 16#01#),
      1732 => to_slv(opcode_type, 16#0A#),
      1733 => to_slv(opcode_type, 16#01#),
      1734 => to_slv(opcode_type, 16#B9#),
      1735 => to_slv(opcode_type, 16#04#),
      1736 => to_slv(opcode_type, 16#01#),
      1737 => to_slv(opcode_type, 16#08#),
      1738 => to_slv(opcode_type, 16#0B#),
      1739 => to_slv(opcode_type, 16#0C#),
      1740 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#09#),
      1761 => to_slv(opcode_type, 16#03#),
      1762 => to_slv(opcode_type, 16#04#),
      1763 => to_slv(opcode_type, 16#08#),
      1764 => to_slv(opcode_type, 16#0D#),
      1765 => to_slv(opcode_type, 16#10#),
      1766 => to_slv(opcode_type, 16#05#),
      1767 => to_slv(opcode_type, 16#07#),
      1768 => to_slv(opcode_type, 16#04#),
      1769 => to_slv(opcode_type, 16#0F#),
      1770 => to_slv(opcode_type, 16#01#),
      1771 => to_slv(opcode_type, 16#0A#),
      1772 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#09#),
      1793 => to_slv(opcode_type, 16#03#),
      1794 => to_slv(opcode_type, 16#01#),
      1795 => to_slv(opcode_type, 16#03#),
      1796 => to_slv(opcode_type, 16#0E#),
      1797 => to_slv(opcode_type, 16#06#),
      1798 => to_slv(opcode_type, 16#03#),
      1799 => to_slv(opcode_type, 16#04#),
      1800 => to_slv(opcode_type, 16#0D#),
      1801 => to_slv(opcode_type, 16#09#),
      1802 => to_slv(opcode_type, 16#0E#),
      1803 => to_slv(opcode_type, 16#0E#),
      1804 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#05#),
      1825 => to_slv(opcode_type, 16#09#),
      1826 => to_slv(opcode_type, 16#02#),
      1827 => to_slv(opcode_type, 16#07#),
      1828 => to_slv(opcode_type, 16#11#),
      1829 => to_slv(opcode_type, 16#0B#),
      1830 => to_slv(opcode_type, 16#08#),
      1831 => to_slv(opcode_type, 16#03#),
      1832 => to_slv(opcode_type, 16#0D#),
      1833 => to_slv(opcode_type, 16#07#),
      1834 => to_slv(opcode_type, 16#0F#),
      1835 => to_slv(opcode_type, 16#0B#),
      1836 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#01#),
      1857 => to_slv(opcode_type, 16#09#),
      1858 => to_slv(opcode_type, 16#07#),
      1859 => to_slv(opcode_type, 16#05#),
      1860 => to_slv(opcode_type, 16#0A#),
      1861 => to_slv(opcode_type, 16#01#),
      1862 => to_slv(opcode_type, 16#0E#),
      1863 => to_slv(opcode_type, 16#08#),
      1864 => to_slv(opcode_type, 16#06#),
      1865 => to_slv(opcode_type, 16#0B#),
      1866 => to_slv(opcode_type, 16#0C#),
      1867 => to_slv(opcode_type, 16#0A#),
      1868 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#07#),
      1890 => to_slv(opcode_type, 16#09#),
      1891 => to_slv(opcode_type, 16#01#),
      1892 => to_slv(opcode_type, 16#80#),
      1893 => to_slv(opcode_type, 16#06#),
      1894 => to_slv(opcode_type, 16#0B#),
      1895 => to_slv(opcode_type, 16#11#),
      1896 => to_slv(opcode_type, 16#06#),
      1897 => to_slv(opcode_type, 16#0F#),
      1898 => to_slv(opcode_type, 16#11#),
      1899 => to_slv(opcode_type, 16#38#),
      1900 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#07#),
      1921 => to_slv(opcode_type, 16#07#),
      1922 => to_slv(opcode_type, 16#08#),
      1923 => to_slv(opcode_type, 16#03#),
      1924 => to_slv(opcode_type, 16#0D#),
      1925 => to_slv(opcode_type, 16#05#),
      1926 => to_slv(opcode_type, 16#0C#),
      1927 => to_slv(opcode_type, 16#07#),
      1928 => to_slv(opcode_type, 16#04#),
      1929 => to_slv(opcode_type, 16#0B#),
      1930 => to_slv(opcode_type, 16#0B#),
      1931 => to_slv(opcode_type, 16#0C#),
      1932 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#08#),
      1953 => to_slv(opcode_type, 16#06#),
      1954 => to_slv(opcode_type, 16#06#),
      1955 => to_slv(opcode_type, 16#09#),
      1956 => to_slv(opcode_type, 16#0A#),
      1957 => to_slv(opcode_type, 16#0E#),
      1958 => to_slv(opcode_type, 16#02#),
      1959 => to_slv(opcode_type, 16#0A#),
      1960 => to_slv(opcode_type, 16#03#),
      1961 => to_slv(opcode_type, 16#05#),
      1962 => to_slv(opcode_type, 16#94#),
      1963 => to_slv(opcode_type, 16#0D#),
      1964 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#07#),
      1985 => to_slv(opcode_type, 16#09#),
      1986 => to_slv(opcode_type, 16#03#),
      1987 => to_slv(opcode_type, 16#09#),
      1988 => to_slv(opcode_type, 16#10#),
      1989 => to_slv(opcode_type, 16#0F#),
      1990 => to_slv(opcode_type, 16#07#),
      1991 => to_slv(opcode_type, 16#08#),
      1992 => to_slv(opcode_type, 16#11#),
      1993 => to_slv(opcode_type, 16#10#),
      1994 => to_slv(opcode_type, 16#11#),
      1995 => to_slv(opcode_type, 16#0D#),
      1996 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#01#),
      2017 => to_slv(opcode_type, 16#07#),
      2018 => to_slv(opcode_type, 16#03#),
      2019 => to_slv(opcode_type, 16#01#),
      2020 => to_slv(opcode_type, 16#10#),
      2021 => to_slv(opcode_type, 16#07#),
      2022 => to_slv(opcode_type, 16#07#),
      2023 => to_slv(opcode_type, 16#10#),
      2024 => to_slv(opcode_type, 16#0A#),
      2025 => to_slv(opcode_type, 16#07#),
      2026 => to_slv(opcode_type, 16#10#),
      2027 => to_slv(opcode_type, 16#0C#),
      2028 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#08#),
      2049 => to_slv(opcode_type, 16#09#),
      2050 => to_slv(opcode_type, 16#08#),
      2051 => to_slv(opcode_type, 16#06#),
      2052 => to_slv(opcode_type, 16#0A#),
      2053 => to_slv(opcode_type, 16#0D#),
      2054 => to_slv(opcode_type, 16#05#),
      2055 => to_slv(opcode_type, 16#0F#),
      2056 => to_slv(opcode_type, 16#08#),
      2057 => to_slv(opcode_type, 16#0B#),
      2058 => to_slv(opcode_type, 16#10#),
      2059 => to_slv(opcode_type, 16#0D#),
      2060 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#03#),
      2081 => to_slv(opcode_type, 16#07#),
      2082 => to_slv(opcode_type, 16#04#),
      2083 => to_slv(opcode_type, 16#09#),
      2084 => to_slv(opcode_type, 16#0E#),
      2085 => to_slv(opcode_type, 16#0A#),
      2086 => to_slv(opcode_type, 16#06#),
      2087 => to_slv(opcode_type, 16#02#),
      2088 => to_slv(opcode_type, 16#0F#),
      2089 => to_slv(opcode_type, 16#09#),
      2090 => to_slv(opcode_type, 16#0B#),
      2091 => to_slv(opcode_type, 16#0C#),
      2092 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#03#),
      2113 => to_slv(opcode_type, 16#09#),
      2114 => to_slv(opcode_type, 16#05#),
      2115 => to_slv(opcode_type, 16#05#),
      2116 => to_slv(opcode_type, 16#3C#),
      2117 => to_slv(opcode_type, 16#09#),
      2118 => to_slv(opcode_type, 16#08#),
      2119 => to_slv(opcode_type, 16#0B#),
      2120 => to_slv(opcode_type, 16#0E#),
      2121 => to_slv(opcode_type, 16#08#),
      2122 => to_slv(opcode_type, 16#0E#),
      2123 => to_slv(opcode_type, 16#0A#),
      2124 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#07#),
      2145 => to_slv(opcode_type, 16#04#),
      2146 => to_slv(opcode_type, 16#06#),
      2147 => to_slv(opcode_type, 16#03#),
      2148 => to_slv(opcode_type, 16#0A#),
      2149 => to_slv(opcode_type, 16#02#),
      2150 => to_slv(opcode_type, 16#0D#),
      2151 => to_slv(opcode_type, 16#04#),
      2152 => to_slv(opcode_type, 16#08#),
      2153 => to_slv(opcode_type, 16#05#),
      2154 => to_slv(opcode_type, 16#11#),
      2155 => to_slv(opcode_type, 16#0A#),
      2156 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#09#),
      2177 => to_slv(opcode_type, 16#09#),
      2178 => to_slv(opcode_type, 16#08#),
      2179 => to_slv(opcode_type, 16#06#),
      2180 => to_slv(opcode_type, 16#0B#),
      2181 => to_slv(opcode_type, 16#0F#),
      2182 => to_slv(opcode_type, 16#08#),
      2183 => to_slv(opcode_type, 16#0D#),
      2184 => to_slv(opcode_type, 16#0F#),
      2185 => to_slv(opcode_type, 16#01#),
      2186 => to_slv(opcode_type, 16#0F#),
      2187 => to_slv(opcode_type, 16#0C#),
      2188 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#06#),
      2209 => to_slv(opcode_type, 16#03#),
      2210 => to_slv(opcode_type, 16#02#),
      2211 => to_slv(opcode_type, 16#04#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#03#),
      2214 => to_slv(opcode_type, 16#08#),
      2215 => to_slv(opcode_type, 16#04#),
      2216 => to_slv(opcode_type, 16#0B#),
      2217 => to_slv(opcode_type, 16#08#),
      2218 => to_slv(opcode_type, 16#0C#),
      2219 => to_slv(opcode_type, 16#0A#),
      2220 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#03#),
      2242 => to_slv(opcode_type, 16#03#),
      2243 => to_slv(opcode_type, 16#09#),
      2244 => to_slv(opcode_type, 16#0F#),
      2245 => to_slv(opcode_type, 16#0E#),
      2246 => to_slv(opcode_type, 16#03#),
      2247 => to_slv(opcode_type, 16#08#),
      2248 => to_slv(opcode_type, 16#08#),
      2249 => to_slv(opcode_type, 16#0B#),
      2250 => to_slv(opcode_type, 16#11#),
      2251 => to_slv(opcode_type, 16#73#),
      2252 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#04#),
      2273 => to_slv(opcode_type, 16#09#),
      2274 => to_slv(opcode_type, 16#09#),
      2275 => to_slv(opcode_type, 16#06#),
      2276 => to_slv(opcode_type, 16#0E#),
      2277 => to_slv(opcode_type, 16#11#),
      2278 => to_slv(opcode_type, 16#04#),
      2279 => to_slv(opcode_type, 16#11#),
      2280 => to_slv(opcode_type, 16#08#),
      2281 => to_slv(opcode_type, 16#03#),
      2282 => to_slv(opcode_type, 16#10#),
      2283 => to_slv(opcode_type, 16#0B#),
      2284 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#02#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#02#),
      2307 => to_slv(opcode_type, 16#01#),
      2308 => to_slv(opcode_type, 16#0D#),
      2309 => to_slv(opcode_type, 16#06#),
      2310 => to_slv(opcode_type, 16#08#),
      2311 => to_slv(opcode_type, 16#0E#),
      2312 => to_slv(opcode_type, 16#0A#),
      2313 => to_slv(opcode_type, 16#08#),
      2314 => to_slv(opcode_type, 16#0A#),
      2315 => to_slv(opcode_type, 16#A9#),
      2316 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#04#),
      2337 => to_slv(opcode_type, 16#08#),
      2338 => to_slv(opcode_type, 16#04#),
      2339 => to_slv(opcode_type, 16#09#),
      2340 => to_slv(opcode_type, 16#10#),
      2341 => to_slv(opcode_type, 16#0D#),
      2342 => to_slv(opcode_type, 16#07#),
      2343 => to_slv(opcode_type, 16#08#),
      2344 => to_slv(opcode_type, 16#11#),
      2345 => to_slv(opcode_type, 16#0E#),
      2346 => to_slv(opcode_type, 16#05#),
      2347 => to_slv(opcode_type, 16#11#),
      2348 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#05#),
      2369 => to_slv(opcode_type, 16#08#),
      2370 => to_slv(opcode_type, 16#05#),
      2371 => to_slv(opcode_type, 16#09#),
      2372 => to_slv(opcode_type, 16#0F#),
      2373 => to_slv(opcode_type, 16#10#),
      2374 => to_slv(opcode_type, 16#09#),
      2375 => to_slv(opcode_type, 16#07#),
      2376 => to_slv(opcode_type, 16#0F#),
      2377 => to_slv(opcode_type, 16#0B#),
      2378 => to_slv(opcode_type, 16#01#),
      2379 => to_slv(opcode_type, 16#0D#),
      2380 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#03#),
      2402 => to_slv(opcode_type, 16#07#),
      2403 => to_slv(opcode_type, 16#01#),
      2404 => to_slv(opcode_type, 16#0E#),
      2405 => to_slv(opcode_type, 16#07#),
      2406 => to_slv(opcode_type, 16#0E#),
      2407 => to_slv(opcode_type, 16#0E#),
      2408 => to_slv(opcode_type, 16#03#),
      2409 => to_slv(opcode_type, 16#01#),
      2410 => to_slv(opcode_type, 16#04#),
      2411 => to_slv(opcode_type, 16#0F#),
      2412 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#09#),
      2433 => to_slv(opcode_type, 16#06#),
      2434 => to_slv(opcode_type, 16#03#),
      2435 => to_slv(opcode_type, 16#01#),
      2436 => to_slv(opcode_type, 16#FD#),
      2437 => to_slv(opcode_type, 16#06#),
      2438 => to_slv(opcode_type, 16#09#),
      2439 => to_slv(opcode_type, 16#0F#),
      2440 => to_slv(opcode_type, 16#0E#),
      2441 => to_slv(opcode_type, 16#02#),
      2442 => to_slv(opcode_type, 16#11#),
      2443 => to_slv(opcode_type, 16#0B#),
      2444 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#09#),
      2465 => to_slv(opcode_type, 16#07#),
      2466 => to_slv(opcode_type, 16#06#),
      2467 => to_slv(opcode_type, 16#04#),
      2468 => to_slv(opcode_type, 16#0C#),
      2469 => to_slv(opcode_type, 16#04#),
      2470 => to_slv(opcode_type, 16#10#),
      2471 => to_slv(opcode_type, 16#08#),
      2472 => to_slv(opcode_type, 16#04#),
      2473 => to_slv(opcode_type, 16#0D#),
      2474 => to_slv(opcode_type, 16#0D#),
      2475 => to_slv(opcode_type, 16#0A#),
      2476 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#01#),
      2497 => to_slv(opcode_type, 16#07#),
      2498 => to_slv(opcode_type, 16#03#),
      2499 => to_slv(opcode_type, 16#05#),
      2500 => to_slv(opcode_type, 16#0E#),
      2501 => to_slv(opcode_type, 16#08#),
      2502 => to_slv(opcode_type, 16#06#),
      2503 => to_slv(opcode_type, 16#10#),
      2504 => to_slv(opcode_type, 16#0C#),
      2505 => to_slv(opcode_type, 16#06#),
      2506 => to_slv(opcode_type, 16#0E#),
      2507 => to_slv(opcode_type, 16#10#),
      2508 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#03#),
      2529 => to_slv(opcode_type, 16#09#),
      2530 => to_slv(opcode_type, 16#06#),
      2531 => to_slv(opcode_type, 16#04#),
      2532 => to_slv(opcode_type, 16#0D#),
      2533 => to_slv(opcode_type, 16#08#),
      2534 => to_slv(opcode_type, 16#11#),
      2535 => to_slv(opcode_type, 16#0D#),
      2536 => to_slv(opcode_type, 16#01#),
      2537 => to_slv(opcode_type, 16#09#),
      2538 => to_slv(opcode_type, 16#0F#),
      2539 => to_slv(opcode_type, 16#10#),
      2540 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#05#),
      2561 => to_slv(opcode_type, 16#09#),
      2562 => to_slv(opcode_type, 16#04#),
      2563 => to_slv(opcode_type, 16#07#),
      2564 => to_slv(opcode_type, 16#0D#),
      2565 => to_slv(opcode_type, 16#0D#),
      2566 => to_slv(opcode_type, 16#07#),
      2567 => to_slv(opcode_type, 16#07#),
      2568 => to_slv(opcode_type, 16#11#),
      2569 => to_slv(opcode_type, 16#0A#),
      2570 => to_slv(opcode_type, 16#01#),
      2571 => to_slv(opcode_type, 16#0B#),
      2572 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#04#),
      2593 => to_slv(opcode_type, 16#06#),
      2594 => to_slv(opcode_type, 16#09#),
      2595 => to_slv(opcode_type, 16#09#),
      2596 => to_slv(opcode_type, 16#0D#),
      2597 => to_slv(opcode_type, 16#0B#),
      2598 => to_slv(opcode_type, 16#09#),
      2599 => to_slv(opcode_type, 16#0D#),
      2600 => to_slv(opcode_type, 16#0F#),
      2601 => to_slv(opcode_type, 16#08#),
      2602 => to_slv(opcode_type, 16#11#),
      2603 => to_slv(opcode_type, 16#0F#),
      2604 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#07#),
      2625 => to_slv(opcode_type, 16#09#),
      2626 => to_slv(opcode_type, 16#07#),
      2627 => to_slv(opcode_type, 16#09#),
      2628 => to_slv(opcode_type, 16#0D#),
      2629 => to_slv(opcode_type, 16#A7#),
      2630 => to_slv(opcode_type, 16#02#),
      2631 => to_slv(opcode_type, 16#0D#),
      2632 => to_slv(opcode_type, 16#02#),
      2633 => to_slv(opcode_type, 16#01#),
      2634 => to_slv(opcode_type, 16#0E#),
      2635 => to_slv(opcode_type, 16#11#),
      2636 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#08#),
      2657 => to_slv(opcode_type, 16#04#),
      2658 => to_slv(opcode_type, 16#09#),
      2659 => to_slv(opcode_type, 16#09#),
      2660 => to_slv(opcode_type, 16#0C#),
      2661 => to_slv(opcode_type, 16#10#),
      2662 => to_slv(opcode_type, 16#09#),
      2663 => to_slv(opcode_type, 16#0E#),
      2664 => to_slv(opcode_type, 16#0C#),
      2665 => to_slv(opcode_type, 16#07#),
      2666 => to_slv(opcode_type, 16#0C#),
      2667 => to_slv(opcode_type, 16#10#),
      2668 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#06#),
      2689 => to_slv(opcode_type, 16#03#),
      2690 => to_slv(opcode_type, 16#07#),
      2691 => to_slv(opcode_type, 16#02#),
      2692 => to_slv(opcode_type, 16#49#),
      2693 => to_slv(opcode_type, 16#03#),
      2694 => to_slv(opcode_type, 16#11#),
      2695 => to_slv(opcode_type, 16#05#),
      2696 => to_slv(opcode_type, 16#08#),
      2697 => to_slv(opcode_type, 16#05#),
      2698 => to_slv(opcode_type, 16#10#),
      2699 => to_slv(opcode_type, 16#10#),
      2700 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#05#),
      2721 => to_slv(opcode_type, 16#08#),
      2722 => to_slv(opcode_type, 16#01#),
      2723 => to_slv(opcode_type, 16#07#),
      2724 => to_slv(opcode_type, 16#0E#),
      2725 => to_slv(opcode_type, 16#11#),
      2726 => to_slv(opcode_type, 16#08#),
      2727 => to_slv(opcode_type, 16#04#),
      2728 => to_slv(opcode_type, 16#0E#),
      2729 => to_slv(opcode_type, 16#08#),
      2730 => to_slv(opcode_type, 16#0D#),
      2731 => to_slv(opcode_type, 16#0A#),
      2732 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#04#),
      2753 => to_slv(opcode_type, 16#06#),
      2754 => to_slv(opcode_type, 16#02#),
      2755 => to_slv(opcode_type, 16#02#),
      2756 => to_slv(opcode_type, 16#0B#),
      2757 => to_slv(opcode_type, 16#06#),
      2758 => to_slv(opcode_type, 16#08#),
      2759 => to_slv(opcode_type, 16#0B#),
      2760 => to_slv(opcode_type, 16#0E#),
      2761 => to_slv(opcode_type, 16#06#),
      2762 => to_slv(opcode_type, 16#0D#),
      2763 => to_slv(opcode_type, 16#10#),
      2764 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#06#),
      2785 => to_slv(opcode_type, 16#02#),
      2786 => to_slv(opcode_type, 16#02#),
      2787 => to_slv(opcode_type, 16#03#),
      2788 => to_slv(opcode_type, 16#0E#),
      2789 => to_slv(opcode_type, 16#03#),
      2790 => to_slv(opcode_type, 16#06#),
      2791 => to_slv(opcode_type, 16#03#),
      2792 => to_slv(opcode_type, 16#0F#),
      2793 => to_slv(opcode_type, 16#06#),
      2794 => to_slv(opcode_type, 16#0E#),
      2795 => to_slv(opcode_type, 16#9D#),
      2796 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#09#),
      2817 => to_slv(opcode_type, 16#04#),
      2818 => to_slv(opcode_type, 16#04#),
      2819 => to_slv(opcode_type, 16#01#),
      2820 => to_slv(opcode_type, 16#10#),
      2821 => to_slv(opcode_type, 16#02#),
      2822 => to_slv(opcode_type, 16#06#),
      2823 => to_slv(opcode_type, 16#08#),
      2824 => to_slv(opcode_type, 16#0B#),
      2825 => to_slv(opcode_type, 16#0D#),
      2826 => to_slv(opcode_type, 16#01#),
      2827 => to_slv(opcode_type, 16#49#),
      2828 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#07#),
      2849 => to_slv(opcode_type, 16#06#),
      2850 => to_slv(opcode_type, 16#01#),
      2851 => to_slv(opcode_type, 16#03#),
      2852 => to_slv(opcode_type, 16#A7#),
      2853 => to_slv(opcode_type, 16#06#),
      2854 => to_slv(opcode_type, 16#02#),
      2855 => to_slv(opcode_type, 16#0D#),
      2856 => to_slv(opcode_type, 16#08#),
      2857 => to_slv(opcode_type, 16#0B#),
      2858 => to_slv(opcode_type, 16#10#),
      2859 => to_slv(opcode_type, 16#0B#),
      2860 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#01#),
      2881 => to_slv(opcode_type, 16#08#),
      2882 => to_slv(opcode_type, 16#02#),
      2883 => to_slv(opcode_type, 16#07#),
      2884 => to_slv(opcode_type, 16#0C#),
      2885 => to_slv(opcode_type, 16#0A#),
      2886 => to_slv(opcode_type, 16#09#),
      2887 => to_slv(opcode_type, 16#08#),
      2888 => to_slv(opcode_type, 16#0D#),
      2889 => to_slv(opcode_type, 16#0C#),
      2890 => to_slv(opcode_type, 16#01#),
      2891 => to_slv(opcode_type, 16#0A#),
      2892 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#07#),
      2913 => to_slv(opcode_type, 16#04#),
      2914 => to_slv(opcode_type, 16#03#),
      2915 => to_slv(opcode_type, 16#01#),
      2916 => to_slv(opcode_type, 16#10#),
      2917 => to_slv(opcode_type, 16#04#),
      2918 => to_slv(opcode_type, 16#09#),
      2919 => to_slv(opcode_type, 16#03#),
      2920 => to_slv(opcode_type, 16#11#),
      2921 => to_slv(opcode_type, 16#08#),
      2922 => to_slv(opcode_type, 16#1E#),
      2923 => to_slv(opcode_type, 16#0D#),
      2924 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#02#),
      2945 => to_slv(opcode_type, 16#08#),
      2946 => to_slv(opcode_type, 16#06#),
      2947 => to_slv(opcode_type, 16#01#),
      2948 => to_slv(opcode_type, 16#0F#),
      2949 => to_slv(opcode_type, 16#07#),
      2950 => to_slv(opcode_type, 16#0C#),
      2951 => to_slv(opcode_type, 16#10#),
      2952 => to_slv(opcode_type, 16#02#),
      2953 => to_slv(opcode_type, 16#08#),
      2954 => to_slv(opcode_type, 16#90#),
      2955 => to_slv(opcode_type, 16#0D#),
      2956 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#05#),
      2977 => to_slv(opcode_type, 16#07#),
      2978 => to_slv(opcode_type, 16#07#),
      2979 => to_slv(opcode_type, 16#03#),
      2980 => to_slv(opcode_type, 16#0C#),
      2981 => to_slv(opcode_type, 16#07#),
      2982 => to_slv(opcode_type, 16#10#),
      2983 => to_slv(opcode_type, 16#0C#),
      2984 => to_slv(opcode_type, 16#02#),
      2985 => to_slv(opcode_type, 16#07#),
      2986 => to_slv(opcode_type, 16#0D#),
      2987 => to_slv(opcode_type, 16#0C#),
      2988 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#04#),
      3009 => to_slv(opcode_type, 16#08#),
      3010 => to_slv(opcode_type, 16#01#),
      3011 => to_slv(opcode_type, 16#02#),
      3012 => to_slv(opcode_type, 16#11#),
      3013 => to_slv(opcode_type, 16#07#),
      3014 => to_slv(opcode_type, 16#06#),
      3015 => to_slv(opcode_type, 16#0F#),
      3016 => to_slv(opcode_type, 16#0F#),
      3017 => to_slv(opcode_type, 16#08#),
      3018 => to_slv(opcode_type, 16#0F#),
      3019 => to_slv(opcode_type, 16#0B#),
      3020 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#02#),
      3041 => to_slv(opcode_type, 16#06#),
      3042 => to_slv(opcode_type, 16#09#),
      3043 => to_slv(opcode_type, 16#05#),
      3044 => to_slv(opcode_type, 16#0B#),
      3045 => to_slv(opcode_type, 16#02#),
      3046 => to_slv(opcode_type, 16#0F#),
      3047 => to_slv(opcode_type, 16#08#),
      3048 => to_slv(opcode_type, 16#01#),
      3049 => to_slv(opcode_type, 16#0B#),
      3050 => to_slv(opcode_type, 16#03#),
      3051 => to_slv(opcode_type, 16#10#),
      3052 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#04#),
      3073 => to_slv(opcode_type, 16#07#),
      3074 => to_slv(opcode_type, 16#07#),
      3075 => to_slv(opcode_type, 16#03#),
      3076 => to_slv(opcode_type, 16#88#),
      3077 => to_slv(opcode_type, 16#07#),
      3078 => to_slv(opcode_type, 16#10#),
      3079 => to_slv(opcode_type, 16#0A#),
      3080 => to_slv(opcode_type, 16#08#),
      3081 => to_slv(opcode_type, 16#03#),
      3082 => to_slv(opcode_type, 16#0D#),
      3083 => to_slv(opcode_type, 16#0E#),
      3084 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#08#),
      3105 => to_slv(opcode_type, 16#09#),
      3106 => to_slv(opcode_type, 16#02#),
      3107 => to_slv(opcode_type, 16#04#),
      3108 => to_slv(opcode_type, 16#0E#),
      3109 => to_slv(opcode_type, 16#05#),
      3110 => to_slv(opcode_type, 16#03#),
      3111 => to_slv(opcode_type, 16#0C#),
      3112 => to_slv(opcode_type, 16#06#),
      3113 => to_slv(opcode_type, 16#02#),
      3114 => to_slv(opcode_type, 16#0A#),
      3115 => to_slv(opcode_type, 16#11#),
      3116 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#05#),
      3137 => to_slv(opcode_type, 16#06#),
      3138 => to_slv(opcode_type, 16#09#),
      3139 => to_slv(opcode_type, 16#01#),
      3140 => to_slv(opcode_type, 16#0C#),
      3141 => to_slv(opcode_type, 16#04#),
      3142 => to_slv(opcode_type, 16#0E#),
      3143 => to_slv(opcode_type, 16#07#),
      3144 => to_slv(opcode_type, 16#09#),
      3145 => to_slv(opcode_type, 16#0D#),
      3146 => to_slv(opcode_type, 16#0F#),
      3147 => to_slv(opcode_type, 16#11#),
      3148 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#04#),
      3169 => to_slv(opcode_type, 16#09#),
      3170 => to_slv(opcode_type, 16#03#),
      3171 => to_slv(opcode_type, 16#02#),
      3172 => to_slv(opcode_type, 16#11#),
      3173 => to_slv(opcode_type, 16#08#),
      3174 => to_slv(opcode_type, 16#09#),
      3175 => to_slv(opcode_type, 16#11#),
      3176 => to_slv(opcode_type, 16#65#),
      3177 => to_slv(opcode_type, 16#06#),
      3178 => to_slv(opcode_type, 16#0D#),
      3179 => to_slv(opcode_type, 16#0B#),
      3180 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#09#),
      3201 => to_slv(opcode_type, 16#08#),
      3202 => to_slv(opcode_type, 16#01#),
      3203 => to_slv(opcode_type, 16#07#),
      3204 => to_slv(opcode_type, 16#0C#),
      3205 => to_slv(opcode_type, 16#0E#),
      3206 => to_slv(opcode_type, 16#07#),
      3207 => to_slv(opcode_type, 16#01#),
      3208 => to_slv(opcode_type, 16#0D#),
      3209 => to_slv(opcode_type, 16#04#),
      3210 => to_slv(opcode_type, 16#11#),
      3211 => to_slv(opcode_type, 16#0F#),
      3212 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#02#),
      3233 => to_slv(opcode_type, 16#08#),
      3234 => to_slv(opcode_type, 16#02#),
      3235 => to_slv(opcode_type, 16#03#),
      3236 => to_slv(opcode_type, 16#11#),
      3237 => to_slv(opcode_type, 16#07#),
      3238 => to_slv(opcode_type, 16#06#),
      3239 => to_slv(opcode_type, 16#0B#),
      3240 => to_slv(opcode_type, 16#0A#),
      3241 => to_slv(opcode_type, 16#09#),
      3242 => to_slv(opcode_type, 16#0B#),
      3243 => to_slv(opcode_type, 16#0D#),
      3244 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#03#),
      3265 => to_slv(opcode_type, 16#07#),
      3266 => to_slv(opcode_type, 16#01#),
      3267 => to_slv(opcode_type, 16#03#),
      3268 => to_slv(opcode_type, 16#0E#),
      3269 => to_slv(opcode_type, 16#06#),
      3270 => to_slv(opcode_type, 16#09#),
      3271 => to_slv(opcode_type, 16#11#),
      3272 => to_slv(opcode_type, 16#0A#),
      3273 => to_slv(opcode_type, 16#07#),
      3274 => to_slv(opcode_type, 16#11#),
      3275 => to_slv(opcode_type, 16#0D#),
      3276 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#02#),
      3297 => to_slv(opcode_type, 16#09#),
      3298 => to_slv(opcode_type, 16#02#),
      3299 => to_slv(opcode_type, 16#05#),
      3300 => to_slv(opcode_type, 16#0E#),
      3301 => to_slv(opcode_type, 16#06#),
      3302 => to_slv(opcode_type, 16#07#),
      3303 => to_slv(opcode_type, 16#0B#),
      3304 => to_slv(opcode_type, 16#51#),
      3305 => to_slv(opcode_type, 16#07#),
      3306 => to_slv(opcode_type, 16#0E#),
      3307 => to_slv(opcode_type, 16#0A#),
      3308 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#07#),
      3329 => to_slv(opcode_type, 16#06#),
      3330 => to_slv(opcode_type, 16#02#),
      3331 => to_slv(opcode_type, 16#02#),
      3332 => to_slv(opcode_type, 16#0B#),
      3333 => to_slv(opcode_type, 16#09#),
      3334 => to_slv(opcode_type, 16#02#),
      3335 => to_slv(opcode_type, 16#10#),
      3336 => to_slv(opcode_type, 16#09#),
      3337 => to_slv(opcode_type, 16#0B#),
      3338 => to_slv(opcode_type, 16#0D#),
      3339 => to_slv(opcode_type, 16#11#),
      3340 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#04#),
      3361 => to_slv(opcode_type, 16#09#),
      3362 => to_slv(opcode_type, 16#08#),
      3363 => to_slv(opcode_type, 16#05#),
      3364 => to_slv(opcode_type, 16#0B#),
      3365 => to_slv(opcode_type, 16#01#),
      3366 => to_slv(opcode_type, 16#11#),
      3367 => to_slv(opcode_type, 16#07#),
      3368 => to_slv(opcode_type, 16#04#),
      3369 => to_slv(opcode_type, 16#10#),
      3370 => to_slv(opcode_type, 16#01#),
      3371 => to_slv(opcode_type, 16#0F#),
      3372 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#09#),
      3393 => to_slv(opcode_type, 16#05#),
      3394 => to_slv(opcode_type, 16#05#),
      3395 => to_slv(opcode_type, 16#02#),
      3396 => to_slv(opcode_type, 16#0C#),
      3397 => to_slv(opcode_type, 16#08#),
      3398 => to_slv(opcode_type, 16#07#),
      3399 => to_slv(opcode_type, 16#03#),
      3400 => to_slv(opcode_type, 16#0D#),
      3401 => to_slv(opcode_type, 16#01#),
      3402 => to_slv(opcode_type, 16#11#),
      3403 => to_slv(opcode_type, 16#0E#),
      3404 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#05#),
      3425 => to_slv(opcode_type, 16#09#),
      3426 => to_slv(opcode_type, 16#08#),
      3427 => to_slv(opcode_type, 16#09#),
      3428 => to_slv(opcode_type, 16#91#),
      3429 => to_slv(opcode_type, 16#10#),
      3430 => to_slv(opcode_type, 16#03#),
      3431 => to_slv(opcode_type, 16#0A#),
      3432 => to_slv(opcode_type, 16#02#),
      3433 => to_slv(opcode_type, 16#06#),
      3434 => to_slv(opcode_type, 16#11#),
      3435 => to_slv(opcode_type, 16#0E#),
      3436 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#09#),
      3457 => to_slv(opcode_type, 16#08#),
      3458 => to_slv(opcode_type, 16#01#),
      3459 => to_slv(opcode_type, 16#06#),
      3460 => to_slv(opcode_type, 16#10#),
      3461 => to_slv(opcode_type, 16#0F#),
      3462 => to_slv(opcode_type, 16#06#),
      3463 => to_slv(opcode_type, 16#02#),
      3464 => to_slv(opcode_type, 16#11#),
      3465 => to_slv(opcode_type, 16#01#),
      3466 => to_slv(opcode_type, 16#0F#),
      3467 => to_slv(opcode_type, 16#0B#),
      3468 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#05#),
      3489 => to_slv(opcode_type, 16#06#),
      3490 => to_slv(opcode_type, 16#06#),
      3491 => to_slv(opcode_type, 16#01#),
      3492 => to_slv(opcode_type, 16#0C#),
      3493 => to_slv(opcode_type, 16#07#),
      3494 => to_slv(opcode_type, 16#0D#),
      3495 => to_slv(opcode_type, 16#10#),
      3496 => to_slv(opcode_type, 16#04#),
      3497 => to_slv(opcode_type, 16#08#),
      3498 => to_slv(opcode_type, 16#0C#),
      3499 => to_slv(opcode_type, 16#0E#),
      3500 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#07#),
      3521 => to_slv(opcode_type, 16#06#),
      3522 => to_slv(opcode_type, 16#05#),
      3523 => to_slv(opcode_type, 16#02#),
      3524 => to_slv(opcode_type, 16#0F#),
      3525 => to_slv(opcode_type, 16#08#),
      3526 => to_slv(opcode_type, 16#08#),
      3527 => to_slv(opcode_type, 16#0F#),
      3528 => to_slv(opcode_type, 16#10#),
      3529 => to_slv(opcode_type, 16#05#),
      3530 => to_slv(opcode_type, 16#0B#),
      3531 => to_slv(opcode_type, 16#10#),
      3532 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#05#),
      3553 => to_slv(opcode_type, 16#07#),
      3554 => to_slv(opcode_type, 16#07#),
      3555 => to_slv(opcode_type, 16#09#),
      3556 => to_slv(opcode_type, 16#0F#),
      3557 => to_slv(opcode_type, 16#0B#),
      3558 => to_slv(opcode_type, 16#01#),
      3559 => to_slv(opcode_type, 16#11#),
      3560 => to_slv(opcode_type, 16#07#),
      3561 => to_slv(opcode_type, 16#02#),
      3562 => to_slv(opcode_type, 16#11#),
      3563 => to_slv(opcode_type, 16#0C#),
      3564 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#02#),
      3585 => to_slv(opcode_type, 16#08#),
      3586 => to_slv(opcode_type, 16#08#),
      3587 => to_slv(opcode_type, 16#07#),
      3588 => to_slv(opcode_type, 16#0C#),
      3589 => to_slv(opcode_type, 16#0B#),
      3590 => to_slv(opcode_type, 16#05#),
      3591 => to_slv(opcode_type, 16#0C#),
      3592 => to_slv(opcode_type, 16#01#),
      3593 => to_slv(opcode_type, 16#07#),
      3594 => to_slv(opcode_type, 16#0B#),
      3595 => to_slv(opcode_type, 16#76#),
      3596 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#07#),
      3617 => to_slv(opcode_type, 16#03#),
      3618 => to_slv(opcode_type, 16#03#),
      3619 => to_slv(opcode_type, 16#04#),
      3620 => to_slv(opcode_type, 16#11#),
      3621 => to_slv(opcode_type, 16#02#),
      3622 => to_slv(opcode_type, 16#09#),
      3623 => to_slv(opcode_type, 16#04#),
      3624 => to_slv(opcode_type, 16#0A#),
      3625 => to_slv(opcode_type, 16#07#),
      3626 => to_slv(opcode_type, 16#11#),
      3627 => to_slv(opcode_type, 16#E9#),
      3628 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#07#),
      3649 => to_slv(opcode_type, 16#06#),
      3650 => to_slv(opcode_type, 16#04#),
      3651 => to_slv(opcode_type, 16#05#),
      3652 => to_slv(opcode_type, 16#0A#),
      3653 => to_slv(opcode_type, 16#07#),
      3654 => to_slv(opcode_type, 16#01#),
      3655 => to_slv(opcode_type, 16#0F#),
      3656 => to_slv(opcode_type, 16#02#),
      3657 => to_slv(opcode_type, 16#11#),
      3658 => to_slv(opcode_type, 16#05#),
      3659 => to_slv(opcode_type, 16#0E#),
      3660 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#01#),
      3681 => to_slv(opcode_type, 16#07#),
      3682 => to_slv(opcode_type, 16#05#),
      3683 => to_slv(opcode_type, 16#08#),
      3684 => to_slv(opcode_type, 16#10#),
      3685 => to_slv(opcode_type, 16#0D#),
      3686 => to_slv(opcode_type, 16#09#),
      3687 => to_slv(opcode_type, 16#06#),
      3688 => to_slv(opcode_type, 16#0D#),
      3689 => to_slv(opcode_type, 16#0F#),
      3690 => to_slv(opcode_type, 16#05#),
      3691 => to_slv(opcode_type, 16#0E#),
      3692 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#01#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#02#),
      3715 => to_slv(opcode_type, 16#02#),
      3716 => to_slv(opcode_type, 16#0A#),
      3717 => to_slv(opcode_type, 16#06#),
      3718 => to_slv(opcode_type, 16#07#),
      3719 => to_slv(opcode_type, 16#0E#),
      3720 => to_slv(opcode_type, 16#10#),
      3721 => to_slv(opcode_type, 16#07#),
      3722 => to_slv(opcode_type, 16#0A#),
      3723 => to_slv(opcode_type, 16#0B#),
      3724 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#01#),
      3745 => to_slv(opcode_type, 16#06#),
      3746 => to_slv(opcode_type, 16#03#),
      3747 => to_slv(opcode_type, 16#02#),
      3748 => to_slv(opcode_type, 16#0A#),
      3749 => to_slv(opcode_type, 16#07#),
      3750 => to_slv(opcode_type, 16#09#),
      3751 => to_slv(opcode_type, 16#0C#),
      3752 => to_slv(opcode_type, 16#0F#),
      3753 => to_slv(opcode_type, 16#07#),
      3754 => to_slv(opcode_type, 16#0C#),
      3755 => to_slv(opcode_type, 16#0E#),
      3756 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#05#),
      3777 => to_slv(opcode_type, 16#06#),
      3778 => to_slv(opcode_type, 16#01#),
      3779 => to_slv(opcode_type, 16#03#),
      3780 => to_slv(opcode_type, 16#10#),
      3781 => to_slv(opcode_type, 16#07#),
      3782 => to_slv(opcode_type, 16#08#),
      3783 => to_slv(opcode_type, 16#0D#),
      3784 => to_slv(opcode_type, 16#10#),
      3785 => to_slv(opcode_type, 16#08#),
      3786 => to_slv(opcode_type, 16#0D#),
      3787 => to_slv(opcode_type, 16#0D#),
      3788 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#05#),
      3809 => to_slv(opcode_type, 16#09#),
      3810 => to_slv(opcode_type, 16#08#),
      3811 => to_slv(opcode_type, 16#02#),
      3812 => to_slv(opcode_type, 16#0D#),
      3813 => to_slv(opcode_type, 16#01#),
      3814 => to_slv(opcode_type, 16#10#),
      3815 => to_slv(opcode_type, 16#08#),
      3816 => to_slv(opcode_type, 16#09#),
      3817 => to_slv(opcode_type, 16#0A#),
      3818 => to_slv(opcode_type, 16#0B#),
      3819 => to_slv(opcode_type, 16#0F#),
      3820 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#09#),
      3841 => to_slv(opcode_type, 16#07#),
      3842 => to_slv(opcode_type, 16#07#),
      3843 => to_slv(opcode_type, 16#03#),
      3844 => to_slv(opcode_type, 16#0F#),
      3845 => to_slv(opcode_type, 16#09#),
      3846 => to_slv(opcode_type, 16#0F#),
      3847 => to_slv(opcode_type, 16#0C#),
      3848 => to_slv(opcode_type, 16#04#),
      3849 => to_slv(opcode_type, 16#05#),
      3850 => to_slv(opcode_type, 16#0F#),
      3851 => to_slv(opcode_type, 16#0B#),
      3852 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#02#),
      3873 => to_slv(opcode_type, 16#08#),
      3874 => to_slv(opcode_type, 16#03#),
      3875 => to_slv(opcode_type, 16#08#),
      3876 => to_slv(opcode_type, 16#10#),
      3877 => to_slv(opcode_type, 16#10#),
      3878 => to_slv(opcode_type, 16#07#),
      3879 => to_slv(opcode_type, 16#01#),
      3880 => to_slv(opcode_type, 16#0A#),
      3881 => to_slv(opcode_type, 16#08#),
      3882 => to_slv(opcode_type, 16#11#),
      3883 => to_slv(opcode_type, 16#0C#),
      3884 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#05#),
      3905 => to_slv(opcode_type, 16#07#),
      3906 => to_slv(opcode_type, 16#06#),
      3907 => to_slv(opcode_type, 16#03#),
      3908 => to_slv(opcode_type, 16#E9#),
      3909 => to_slv(opcode_type, 16#08#),
      3910 => to_slv(opcode_type, 16#0C#),
      3911 => to_slv(opcode_type, 16#0D#),
      3912 => to_slv(opcode_type, 16#08#),
      3913 => to_slv(opcode_type, 16#03#),
      3914 => to_slv(opcode_type, 16#0C#),
      3915 => to_slv(opcode_type, 16#0A#),
      3916 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#03#),
      3937 => to_slv(opcode_type, 16#09#),
      3938 => to_slv(opcode_type, 16#06#),
      3939 => to_slv(opcode_type, 16#06#),
      3940 => to_slv(opcode_type, 16#C7#),
      3941 => to_slv(opcode_type, 16#0B#),
      3942 => to_slv(opcode_type, 16#07#),
      3943 => to_slv(opcode_type, 16#10#),
      3944 => to_slv(opcode_type, 16#52#),
      3945 => to_slv(opcode_type, 16#03#),
      3946 => to_slv(opcode_type, 16#04#),
      3947 => to_slv(opcode_type, 16#0C#),
      3948 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#03#),
      3969 => to_slv(opcode_type, 16#08#),
      3970 => to_slv(opcode_type, 16#06#),
      3971 => to_slv(opcode_type, 16#09#),
      3972 => to_slv(opcode_type, 16#0B#),
      3973 => to_slv(opcode_type, 16#0C#),
      3974 => to_slv(opcode_type, 16#03#),
      3975 => to_slv(opcode_type, 16#0F#),
      3976 => to_slv(opcode_type, 16#07#),
      3977 => to_slv(opcode_type, 16#05#),
      3978 => to_slv(opcode_type, 16#0C#),
      3979 => to_slv(opcode_type, 16#11#),
      3980 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#05#),
      4001 => to_slv(opcode_type, 16#09#),
      4002 => to_slv(opcode_type, 16#05#),
      4003 => to_slv(opcode_type, 16#09#),
      4004 => to_slv(opcode_type, 16#0E#),
      4005 => to_slv(opcode_type, 16#0E#),
      4006 => to_slv(opcode_type, 16#06#),
      4007 => to_slv(opcode_type, 16#04#),
      4008 => to_slv(opcode_type, 16#0A#),
      4009 => to_slv(opcode_type, 16#09#),
      4010 => to_slv(opcode_type, 16#0F#),
      4011 => to_slv(opcode_type, 16#0E#),
      4012 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#07#),
      4033 => to_slv(opcode_type, 16#08#),
      4034 => to_slv(opcode_type, 16#03#),
      4035 => to_slv(opcode_type, 16#06#),
      4036 => to_slv(opcode_type, 16#5B#),
      4037 => to_slv(opcode_type, 16#0D#),
      4038 => to_slv(opcode_type, 16#08#),
      4039 => to_slv(opcode_type, 16#09#),
      4040 => to_slv(opcode_type, 16#0B#),
      4041 => to_slv(opcode_type, 16#4E#),
      4042 => to_slv(opcode_type, 16#0D#),
      4043 => to_slv(opcode_type, 16#0C#),
      4044 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#07#),
      4065 => to_slv(opcode_type, 16#02#),
      4066 => to_slv(opcode_type, 16#06#),
      4067 => to_slv(opcode_type, 16#05#),
      4068 => to_slv(opcode_type, 16#17#),
      4069 => to_slv(opcode_type, 16#07#),
      4070 => to_slv(opcode_type, 16#0D#),
      4071 => to_slv(opcode_type, 16#0E#),
      4072 => to_slv(opcode_type, 16#04#),
      4073 => to_slv(opcode_type, 16#04#),
      4074 => to_slv(opcode_type, 16#02#),
      4075 => to_slv(opcode_type, 16#8D#),
      4076 to 4095 => (others => '0')
  ),

    -- Bin `13`...
    12 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#08#),
      1 => to_slv(opcode_type, 16#03#),
      2 => to_slv(opcode_type, 16#05#),
      3 => to_slv(opcode_type, 16#01#),
      4 => to_slv(opcode_type, 16#0D#),
      5 => to_slv(opcode_type, 16#04#),
      6 => to_slv(opcode_type, 16#06#),
      7 => to_slv(opcode_type, 16#08#),
      8 => to_slv(opcode_type, 16#10#),
      9 => to_slv(opcode_type, 16#0F#),
      10 => to_slv(opcode_type, 16#06#),
      11 => to_slv(opcode_type, 16#0E#),
      12 => to_slv(opcode_type, 16#C7#),
      13 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#09#),
      33 => to_slv(opcode_type, 16#04#),
      34 => to_slv(opcode_type, 16#01#),
      35 => to_slv(opcode_type, 16#03#),
      36 => to_slv(opcode_type, 16#11#),
      37 => to_slv(opcode_type, 16#01#),
      38 => to_slv(opcode_type, 16#09#),
      39 => to_slv(opcode_type, 16#08#),
      40 => to_slv(opcode_type, 16#0F#),
      41 => to_slv(opcode_type, 16#11#),
      42 => to_slv(opcode_type, 16#07#),
      43 => to_slv(opcode_type, 16#32#),
      44 => to_slv(opcode_type, 16#0A#),
      45 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#05#),
      65 => to_slv(opcode_type, 16#09#),
      66 => to_slv(opcode_type, 16#03#),
      67 => to_slv(opcode_type, 16#07#),
      68 => to_slv(opcode_type, 16#0B#),
      69 => to_slv(opcode_type, 16#0F#),
      70 => to_slv(opcode_type, 16#08#),
      71 => to_slv(opcode_type, 16#09#),
      72 => to_slv(opcode_type, 16#0D#),
      73 => to_slv(opcode_type, 16#0C#),
      74 => to_slv(opcode_type, 16#08#),
      75 => to_slv(opcode_type, 16#0E#),
      76 => to_slv(opcode_type, 16#0D#),
      77 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#08#),
      97 => to_slv(opcode_type, 16#01#),
      98 => to_slv(opcode_type, 16#01#),
      99 => to_slv(opcode_type, 16#09#),
      100 => to_slv(opcode_type, 16#0F#),
      101 => to_slv(opcode_type, 16#C7#),
      102 => to_slv(opcode_type, 16#08#),
      103 => to_slv(opcode_type, 16#07#),
      104 => to_slv(opcode_type, 16#05#),
      105 => to_slv(opcode_type, 16#0E#),
      106 => to_slv(opcode_type, 16#01#),
      107 => to_slv(opcode_type, 16#11#),
      108 => to_slv(opcode_type, 16#10#),
      109 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#08#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#01#),
      131 => to_slv(opcode_type, 16#08#),
      132 => to_slv(opcode_type, 16#0E#),
      133 => to_slv(opcode_type, 16#0F#),
      134 => to_slv(opcode_type, 16#06#),
      135 => to_slv(opcode_type, 16#09#),
      136 => to_slv(opcode_type, 16#0E#),
      137 => to_slv(opcode_type, 16#DE#),
      138 => to_slv(opcode_type, 16#01#),
      139 => to_slv(opcode_type, 16#0C#),
      140 => to_slv(opcode_type, 16#0E#),
      141 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#05#),
      161 => to_slv(opcode_type, 16#08#),
      162 => to_slv(opcode_type, 16#03#),
      163 => to_slv(opcode_type, 16#06#),
      164 => to_slv(opcode_type, 16#D9#),
      165 => to_slv(opcode_type, 16#11#),
      166 => to_slv(opcode_type, 16#09#),
      167 => to_slv(opcode_type, 16#08#),
      168 => to_slv(opcode_type, 16#0D#),
      169 => to_slv(opcode_type, 16#0D#),
      170 => to_slv(opcode_type, 16#09#),
      171 => to_slv(opcode_type, 16#11#),
      172 => to_slv(opcode_type, 16#0A#),
      173 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#01#),
      193 => to_slv(opcode_type, 16#07#),
      194 => to_slv(opcode_type, 16#03#),
      195 => to_slv(opcode_type, 16#06#),
      196 => to_slv(opcode_type, 16#0C#),
      197 => to_slv(opcode_type, 16#0B#),
      198 => to_slv(opcode_type, 16#08#),
      199 => to_slv(opcode_type, 16#08#),
      200 => to_slv(opcode_type, 16#0A#),
      201 => to_slv(opcode_type, 16#0F#),
      202 => to_slv(opcode_type, 16#08#),
      203 => to_slv(opcode_type, 16#0E#),
      204 => to_slv(opcode_type, 16#0C#),
      205 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#08#),
      225 => to_slv(opcode_type, 16#08#),
      226 => to_slv(opcode_type, 16#03#),
      227 => to_slv(opcode_type, 16#04#),
      228 => to_slv(opcode_type, 16#0F#),
      229 => to_slv(opcode_type, 16#08#),
      230 => to_slv(opcode_type, 16#04#),
      231 => to_slv(opcode_type, 16#11#),
      232 => to_slv(opcode_type, 16#05#),
      233 => to_slv(opcode_type, 16#0F#),
      234 => to_slv(opcode_type, 16#07#),
      235 => to_slv(opcode_type, 16#10#),
      236 => to_slv(opcode_type, 16#0E#),
      237 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#07#),
      257 => to_slv(opcode_type, 16#01#),
      258 => to_slv(opcode_type, 16#06#),
      259 => to_slv(opcode_type, 16#07#),
      260 => to_slv(opcode_type, 16#11#),
      261 => to_slv(opcode_type, 16#3D#),
      262 => to_slv(opcode_type, 16#06#),
      263 => to_slv(opcode_type, 16#0C#),
      264 => to_slv(opcode_type, 16#0D#),
      265 => to_slv(opcode_type, 16#06#),
      266 => to_slv(opcode_type, 16#02#),
      267 => to_slv(opcode_type, 16#10#),
      268 => to_slv(opcode_type, 16#0D#),
      269 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#01#),
      289 => to_slv(opcode_type, 16#06#),
      290 => to_slv(opcode_type, 16#09#),
      291 => to_slv(opcode_type, 16#02#),
      292 => to_slv(opcode_type, 16#0C#),
      293 => to_slv(opcode_type, 16#05#),
      294 => to_slv(opcode_type, 16#FF#),
      295 => to_slv(opcode_type, 16#07#),
      296 => to_slv(opcode_type, 16#07#),
      297 => to_slv(opcode_type, 16#0D#),
      298 => to_slv(opcode_type, 16#10#),
      299 => to_slv(opcode_type, 16#02#),
      300 => to_slv(opcode_type, 16#54#),
      301 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#04#),
      321 => to_slv(opcode_type, 16#06#),
      322 => to_slv(opcode_type, 16#05#),
      323 => to_slv(opcode_type, 16#08#),
      324 => to_slv(opcode_type, 16#0B#),
      325 => to_slv(opcode_type, 16#11#),
      326 => to_slv(opcode_type, 16#09#),
      327 => to_slv(opcode_type, 16#09#),
      328 => to_slv(opcode_type, 16#11#),
      329 => to_slv(opcode_type, 16#0C#),
      330 => to_slv(opcode_type, 16#09#),
      331 => to_slv(opcode_type, 16#0C#),
      332 => to_slv(opcode_type, 16#10#),
      333 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#04#),
      353 => to_slv(opcode_type, 16#06#),
      354 => to_slv(opcode_type, 16#07#),
      355 => to_slv(opcode_type, 16#07#),
      356 => to_slv(opcode_type, 16#0B#),
      357 => to_slv(opcode_type, 16#B0#),
      358 => to_slv(opcode_type, 16#08#),
      359 => to_slv(opcode_type, 16#B7#),
      360 => to_slv(opcode_type, 16#0B#),
      361 => to_slv(opcode_type, 16#06#),
      362 => to_slv(opcode_type, 16#01#),
      363 => to_slv(opcode_type, 16#11#),
      364 => to_slv(opcode_type, 16#0F#),
      365 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#02#),
      385 => to_slv(opcode_type, 16#09#),
      386 => to_slv(opcode_type, 16#01#),
      387 => to_slv(opcode_type, 16#09#),
      388 => to_slv(opcode_type, 16#0F#),
      389 => to_slv(opcode_type, 16#0E#),
      390 => to_slv(opcode_type, 16#06#),
      391 => to_slv(opcode_type, 16#08#),
      392 => to_slv(opcode_type, 16#0A#),
      393 => to_slv(opcode_type, 16#3A#),
      394 => to_slv(opcode_type, 16#06#),
      395 => to_slv(opcode_type, 16#10#),
      396 => to_slv(opcode_type, 16#0D#),
      397 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#05#),
      417 => to_slv(opcode_type, 16#06#),
      418 => to_slv(opcode_type, 16#01#),
      419 => to_slv(opcode_type, 16#09#),
      420 => to_slv(opcode_type, 16#0A#),
      421 => to_slv(opcode_type, 16#11#),
      422 => to_slv(opcode_type, 16#07#),
      423 => to_slv(opcode_type, 16#06#),
      424 => to_slv(opcode_type, 16#10#),
      425 => to_slv(opcode_type, 16#59#),
      426 => to_slv(opcode_type, 16#07#),
      427 => to_slv(opcode_type, 16#0F#),
      428 => to_slv(opcode_type, 16#0A#),
      429 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#04#),
      449 => to_slv(opcode_type, 16#08#),
      450 => to_slv(opcode_type, 16#03#),
      451 => to_slv(opcode_type, 16#08#),
      452 => to_slv(opcode_type, 16#0A#),
      453 => to_slv(opcode_type, 16#11#),
      454 => to_slv(opcode_type, 16#06#),
      455 => to_slv(opcode_type, 16#09#),
      456 => to_slv(opcode_type, 16#0A#),
      457 => to_slv(opcode_type, 16#0D#),
      458 => to_slv(opcode_type, 16#08#),
      459 => to_slv(opcode_type, 16#10#),
      460 => to_slv(opcode_type, 16#0A#),
      461 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#09#),
      481 => to_slv(opcode_type, 16#04#),
      482 => to_slv(opcode_type, 16#01#),
      483 => to_slv(opcode_type, 16#08#),
      484 => to_slv(opcode_type, 16#79#),
      485 => to_slv(opcode_type, 16#0B#),
      486 => to_slv(opcode_type, 16#08#),
      487 => to_slv(opcode_type, 16#08#),
      488 => to_slv(opcode_type, 16#03#),
      489 => to_slv(opcode_type, 16#0C#),
      490 => to_slv(opcode_type, 16#01#),
      491 => to_slv(opcode_type, 16#11#),
      492 => to_slv(opcode_type, 16#10#),
      493 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#02#),
      513 => to_slv(opcode_type, 16#08#),
      514 => to_slv(opcode_type, 16#06#),
      515 => to_slv(opcode_type, 16#08#),
      516 => to_slv(opcode_type, 16#0B#),
      517 => to_slv(opcode_type, 16#0E#),
      518 => to_slv(opcode_type, 16#08#),
      519 => to_slv(opcode_type, 16#0B#),
      520 => to_slv(opcode_type, 16#97#),
      521 => to_slv(opcode_type, 16#02#),
      522 => to_slv(opcode_type, 16#09#),
      523 => to_slv(opcode_type, 16#0D#),
      524 => to_slv(opcode_type, 16#0F#),
      525 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#08#),
      545 => to_slv(opcode_type, 16#06#),
      546 => to_slv(opcode_type, 16#05#),
      547 => to_slv(opcode_type, 16#01#),
      548 => to_slv(opcode_type, 16#4B#),
      549 => to_slv(opcode_type, 16#07#),
      550 => to_slv(opcode_type, 16#07#),
      551 => to_slv(opcode_type, 16#9B#),
      552 => to_slv(opcode_type, 16#0D#),
      553 => to_slv(opcode_type, 16#09#),
      554 => to_slv(opcode_type, 16#0E#),
      555 => to_slv(opcode_type, 16#0E#),
      556 => to_slv(opcode_type, 16#5C#),
      557 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#07#),
      577 => to_slv(opcode_type, 16#09#),
      578 => to_slv(opcode_type, 16#02#),
      579 => to_slv(opcode_type, 16#06#),
      580 => to_slv(opcode_type, 16#0C#),
      581 => to_slv(opcode_type, 16#0A#),
      582 => to_slv(opcode_type, 16#04#),
      583 => to_slv(opcode_type, 16#07#),
      584 => to_slv(opcode_type, 16#0F#),
      585 => to_slv(opcode_type, 16#0F#),
      586 => to_slv(opcode_type, 16#07#),
      587 => to_slv(opcode_type, 16#30#),
      588 => to_slv(opcode_type, 16#0E#),
      589 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#04#),
      609 => to_slv(opcode_type, 16#08#),
      610 => to_slv(opcode_type, 16#02#),
      611 => to_slv(opcode_type, 16#07#),
      612 => to_slv(opcode_type, 16#0A#),
      613 => to_slv(opcode_type, 16#D2#),
      614 => to_slv(opcode_type, 16#09#),
      615 => to_slv(opcode_type, 16#07#),
      616 => to_slv(opcode_type, 16#7C#),
      617 => to_slv(opcode_type, 16#0B#),
      618 => to_slv(opcode_type, 16#09#),
      619 => to_slv(opcode_type, 16#11#),
      620 => to_slv(opcode_type, 16#5C#),
      621 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#01#),
      641 => to_slv(opcode_type, 16#08#),
      642 => to_slv(opcode_type, 16#05#),
      643 => to_slv(opcode_type, 16#06#),
      644 => to_slv(opcode_type, 16#0F#),
      645 => to_slv(opcode_type, 16#51#),
      646 => to_slv(opcode_type, 16#09#),
      647 => to_slv(opcode_type, 16#08#),
      648 => to_slv(opcode_type, 16#1E#),
      649 => to_slv(opcode_type, 16#11#),
      650 => to_slv(opcode_type, 16#06#),
      651 => to_slv(opcode_type, 16#0B#),
      652 => to_slv(opcode_type, 16#0E#),
      653 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#04#),
      673 => to_slv(opcode_type, 16#06#),
      674 => to_slv(opcode_type, 16#02#),
      675 => to_slv(opcode_type, 16#07#),
      676 => to_slv(opcode_type, 16#0C#),
      677 => to_slv(opcode_type, 16#10#),
      678 => to_slv(opcode_type, 16#08#),
      679 => to_slv(opcode_type, 16#09#),
      680 => to_slv(opcode_type, 16#0A#),
      681 => to_slv(opcode_type, 16#0A#),
      682 => to_slv(opcode_type, 16#06#),
      683 => to_slv(opcode_type, 16#0D#),
      684 => to_slv(opcode_type, 16#0B#),
      685 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#07#),
      705 => to_slv(opcode_type, 16#03#),
      706 => to_slv(opcode_type, 16#05#),
      707 => to_slv(opcode_type, 16#01#),
      708 => to_slv(opcode_type, 16#0F#),
      709 => to_slv(opcode_type, 16#07#),
      710 => to_slv(opcode_type, 16#05#),
      711 => to_slv(opcode_type, 16#09#),
      712 => to_slv(opcode_type, 16#0B#),
      713 => to_slv(opcode_type, 16#0A#),
      714 => to_slv(opcode_type, 16#08#),
      715 => to_slv(opcode_type, 16#0D#),
      716 => to_slv(opcode_type, 16#0C#),
      717 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#08#),
      737 => to_slv(opcode_type, 16#01#),
      738 => to_slv(opcode_type, 16#02#),
      739 => to_slv(opcode_type, 16#05#),
      740 => to_slv(opcode_type, 16#0E#),
      741 => to_slv(opcode_type, 16#03#),
      742 => to_slv(opcode_type, 16#06#),
      743 => to_slv(opcode_type, 16#07#),
      744 => to_slv(opcode_type, 16#0A#),
      745 => to_slv(opcode_type, 16#0F#),
      746 => to_slv(opcode_type, 16#07#),
      747 => to_slv(opcode_type, 16#4B#),
      748 => to_slv(opcode_type, 16#0B#),
      749 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#06#),
      769 => to_slv(opcode_type, 16#05#),
      770 => to_slv(opcode_type, 16#09#),
      771 => to_slv(opcode_type, 16#04#),
      772 => to_slv(opcode_type, 16#10#),
      773 => to_slv(opcode_type, 16#05#),
      774 => to_slv(opcode_type, 16#10#),
      775 => to_slv(opcode_type, 16#08#),
      776 => to_slv(opcode_type, 16#01#),
      777 => to_slv(opcode_type, 16#05#),
      778 => to_slv(opcode_type, 16#0B#),
      779 => to_slv(opcode_type, 16#05#),
      780 => to_slv(opcode_type, 16#0F#),
      781 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#06#),
      801 => to_slv(opcode_type, 16#09#),
      802 => to_slv(opcode_type, 16#04#),
      803 => to_slv(opcode_type, 16#05#),
      804 => to_slv(opcode_type, 16#0F#),
      805 => to_slv(opcode_type, 16#04#),
      806 => to_slv(opcode_type, 16#03#),
      807 => to_slv(opcode_type, 16#0D#),
      808 => to_slv(opcode_type, 16#04#),
      809 => to_slv(opcode_type, 16#07#),
      810 => to_slv(opcode_type, 16#04#),
      811 => to_slv(opcode_type, 16#11#),
      812 => to_slv(opcode_type, 16#0E#),
      813 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#01#),
      833 => to_slv(opcode_type, 16#06#),
      834 => to_slv(opcode_type, 16#05#),
      835 => to_slv(opcode_type, 16#09#),
      836 => to_slv(opcode_type, 16#0B#),
      837 => to_slv(opcode_type, 16#0A#),
      838 => to_slv(opcode_type, 16#09#),
      839 => to_slv(opcode_type, 16#06#),
      840 => to_slv(opcode_type, 16#11#),
      841 => to_slv(opcode_type, 16#0B#),
      842 => to_slv(opcode_type, 16#07#),
      843 => to_slv(opcode_type, 16#11#),
      844 => to_slv(opcode_type, 16#0D#),
      845 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#06#),
      865 => to_slv(opcode_type, 16#01#),
      866 => to_slv(opcode_type, 16#03#),
      867 => to_slv(opcode_type, 16#09#),
      868 => to_slv(opcode_type, 16#0F#),
      869 => to_slv(opcode_type, 16#10#),
      870 => to_slv(opcode_type, 16#04#),
      871 => to_slv(opcode_type, 16#06#),
      872 => to_slv(opcode_type, 16#08#),
      873 => to_slv(opcode_type, 16#11#),
      874 => to_slv(opcode_type, 16#0A#),
      875 => to_slv(opcode_type, 16#01#),
      876 => to_slv(opcode_type, 16#11#),
      877 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#03#),
      897 => to_slv(opcode_type, 16#08#),
      898 => to_slv(opcode_type, 16#09#),
      899 => to_slv(opcode_type, 16#06#),
      900 => to_slv(opcode_type, 16#0E#),
      901 => to_slv(opcode_type, 16#3D#),
      902 => to_slv(opcode_type, 16#09#),
      903 => to_slv(opcode_type, 16#11#),
      904 => to_slv(opcode_type, 16#0B#),
      905 => to_slv(opcode_type, 16#02#),
      906 => to_slv(opcode_type, 16#09#),
      907 => to_slv(opcode_type, 16#0E#),
      908 => to_slv(opcode_type, 16#10#),
      909 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#01#),
      929 => to_slv(opcode_type, 16#08#),
      930 => to_slv(opcode_type, 16#05#),
      931 => to_slv(opcode_type, 16#06#),
      932 => to_slv(opcode_type, 16#0B#),
      933 => to_slv(opcode_type, 16#0A#),
      934 => to_slv(opcode_type, 16#08#),
      935 => to_slv(opcode_type, 16#08#),
      936 => to_slv(opcode_type, 16#0C#),
      937 => to_slv(opcode_type, 16#19#),
      938 => to_slv(opcode_type, 16#06#),
      939 => to_slv(opcode_type, 16#10#),
      940 => to_slv(opcode_type, 16#10#),
      941 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#04#),
      961 => to_slv(opcode_type, 16#09#),
      962 => to_slv(opcode_type, 16#04#),
      963 => to_slv(opcode_type, 16#09#),
      964 => to_slv(opcode_type, 16#0C#),
      965 => to_slv(opcode_type, 16#0D#),
      966 => to_slv(opcode_type, 16#09#),
      967 => to_slv(opcode_type, 16#06#),
      968 => to_slv(opcode_type, 16#0A#),
      969 => to_slv(opcode_type, 16#A9#),
      970 => to_slv(opcode_type, 16#08#),
      971 => to_slv(opcode_type, 16#0F#),
      972 => to_slv(opcode_type, 16#11#),
      973 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#01#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#06#),
      995 => to_slv(opcode_type, 16#03#),
      996 => to_slv(opcode_type, 16#0A#),
      997 => to_slv(opcode_type, 16#07#),
      998 => to_slv(opcode_type, 16#10#),
      999 => to_slv(opcode_type, 16#11#),
      1000 => to_slv(opcode_type, 16#06#),
      1001 => to_slv(opcode_type, 16#07#),
      1002 => to_slv(opcode_type, 16#10#),
      1003 => to_slv(opcode_type, 16#0D#),
      1004 => to_slv(opcode_type, 16#10#),
      1005 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#06#),
      1025 => to_slv(opcode_type, 16#03#),
      1026 => to_slv(opcode_type, 16#03#),
      1027 => to_slv(opcode_type, 16#08#),
      1028 => to_slv(opcode_type, 16#0A#),
      1029 => to_slv(opcode_type, 16#0C#),
      1030 => to_slv(opcode_type, 16#08#),
      1031 => to_slv(opcode_type, 16#07#),
      1032 => to_slv(opcode_type, 16#05#),
      1033 => to_slv(opcode_type, 16#28#),
      1034 => to_slv(opcode_type, 16#05#),
      1035 => to_slv(opcode_type, 16#0E#),
      1036 => to_slv(opcode_type, 16#0B#),
      1037 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#06#),
      1057 => to_slv(opcode_type, 16#06#),
      1058 => to_slv(opcode_type, 16#08#),
      1059 => to_slv(opcode_type, 16#03#),
      1060 => to_slv(opcode_type, 16#0B#),
      1061 => to_slv(opcode_type, 16#04#),
      1062 => to_slv(opcode_type, 16#0F#),
      1063 => to_slv(opcode_type, 16#09#),
      1064 => to_slv(opcode_type, 16#06#),
      1065 => to_slv(opcode_type, 16#0D#),
      1066 => to_slv(opcode_type, 16#0C#),
      1067 => to_slv(opcode_type, 16#0A#),
      1068 => to_slv(opcode_type, 16#10#),
      1069 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#07#),
      1089 => to_slv(opcode_type, 16#08#),
      1090 => to_slv(opcode_type, 16#04#),
      1091 => to_slv(opcode_type, 16#02#),
      1092 => to_slv(opcode_type, 16#11#),
      1093 => to_slv(opcode_type, 16#03#),
      1094 => to_slv(opcode_type, 16#07#),
      1095 => to_slv(opcode_type, 16#11#),
      1096 => to_slv(opcode_type, 16#0F#),
      1097 => to_slv(opcode_type, 16#04#),
      1098 => to_slv(opcode_type, 16#07#),
      1099 => to_slv(opcode_type, 16#0E#),
      1100 => to_slv(opcode_type, 16#0B#),
      1101 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#09#),
      1121 => to_slv(opcode_type, 16#06#),
      1122 => to_slv(opcode_type, 16#02#),
      1123 => to_slv(opcode_type, 16#06#),
      1124 => to_slv(opcode_type, 16#0D#),
      1125 => to_slv(opcode_type, 16#0E#),
      1126 => to_slv(opcode_type, 16#05#),
      1127 => to_slv(opcode_type, 16#02#),
      1128 => to_slv(opcode_type, 16#0E#),
      1129 => to_slv(opcode_type, 16#07#),
      1130 => to_slv(opcode_type, 16#01#),
      1131 => to_slv(opcode_type, 16#10#),
      1132 => to_slv(opcode_type, 16#0C#),
      1133 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#08#),
      1153 => to_slv(opcode_type, 16#01#),
      1154 => to_slv(opcode_type, 16#09#),
      1155 => to_slv(opcode_type, 16#06#),
      1156 => to_slv(opcode_type, 16#0C#),
      1157 => to_slv(opcode_type, 16#0A#),
      1158 => to_slv(opcode_type, 16#04#),
      1159 => to_slv(opcode_type, 16#DF#),
      1160 => to_slv(opcode_type, 16#03#),
      1161 => to_slv(opcode_type, 16#06#),
      1162 => to_slv(opcode_type, 16#01#),
      1163 => to_slv(opcode_type, 16#B2#),
      1164 => to_slv(opcode_type, 16#0E#),
      1165 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#03#),
      1185 => to_slv(opcode_type, 16#06#),
      1186 => to_slv(opcode_type, 16#07#),
      1187 => to_slv(opcode_type, 16#02#),
      1188 => to_slv(opcode_type, 16#78#),
      1189 => to_slv(opcode_type, 16#06#),
      1190 => to_slv(opcode_type, 16#0A#),
      1191 => to_slv(opcode_type, 16#0A#),
      1192 => to_slv(opcode_type, 16#07#),
      1193 => to_slv(opcode_type, 16#07#),
      1194 => to_slv(opcode_type, 16#0D#),
      1195 => to_slv(opcode_type, 16#0E#),
      1196 => to_slv(opcode_type, 16#0D#),
      1197 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#04#),
      1217 => to_slv(opcode_type, 16#08#),
      1218 => to_slv(opcode_type, 16#05#),
      1219 => to_slv(opcode_type, 16#09#),
      1220 => to_slv(opcode_type, 16#0B#),
      1221 => to_slv(opcode_type, 16#10#),
      1222 => to_slv(opcode_type, 16#08#),
      1223 => to_slv(opcode_type, 16#08#),
      1224 => to_slv(opcode_type, 16#C8#),
      1225 => to_slv(opcode_type, 16#0D#),
      1226 => to_slv(opcode_type, 16#06#),
      1227 => to_slv(opcode_type, 16#0D#),
      1228 => to_slv(opcode_type, 16#0B#),
      1229 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#04#),
      1249 => to_slv(opcode_type, 16#08#),
      1250 => to_slv(opcode_type, 16#09#),
      1251 => to_slv(opcode_type, 16#08#),
      1252 => to_slv(opcode_type, 16#84#),
      1253 => to_slv(opcode_type, 16#0F#),
      1254 => to_slv(opcode_type, 16#03#),
      1255 => to_slv(opcode_type, 16#0E#),
      1256 => to_slv(opcode_type, 16#08#),
      1257 => to_slv(opcode_type, 16#01#),
      1258 => to_slv(opcode_type, 16#10#),
      1259 => to_slv(opcode_type, 16#02#),
      1260 => to_slv(opcode_type, 16#10#),
      1261 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#06#),
      1281 => to_slv(opcode_type, 16#03#),
      1282 => to_slv(opcode_type, 16#07#),
      1283 => to_slv(opcode_type, 16#09#),
      1284 => to_slv(opcode_type, 16#10#),
      1285 => to_slv(opcode_type, 16#3E#),
      1286 => to_slv(opcode_type, 16#04#),
      1287 => to_slv(opcode_type, 16#F4#),
      1288 => to_slv(opcode_type, 16#09#),
      1289 => to_slv(opcode_type, 16#07#),
      1290 => to_slv(opcode_type, 16#0F#),
      1291 => to_slv(opcode_type, 16#0B#),
      1292 => to_slv(opcode_type, 16#0D#),
      1293 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#07#),
      1313 => to_slv(opcode_type, 16#05#),
      1314 => to_slv(opcode_type, 16#08#),
      1315 => to_slv(opcode_type, 16#09#),
      1316 => to_slv(opcode_type, 16#D4#),
      1317 => to_slv(opcode_type, 16#0A#),
      1318 => to_slv(opcode_type, 16#09#),
      1319 => to_slv(opcode_type, 16#0C#),
      1320 => to_slv(opcode_type, 16#11#),
      1321 => to_slv(opcode_type, 16#07#),
      1322 => to_slv(opcode_type, 16#02#),
      1323 => to_slv(opcode_type, 16#0E#),
      1324 => to_slv(opcode_type, 16#10#),
      1325 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#02#),
      1345 => to_slv(opcode_type, 16#08#),
      1346 => to_slv(opcode_type, 16#04#),
      1347 => to_slv(opcode_type, 16#09#),
      1348 => to_slv(opcode_type, 16#10#),
      1349 => to_slv(opcode_type, 16#0A#),
      1350 => to_slv(opcode_type, 16#09#),
      1351 => to_slv(opcode_type, 16#09#),
      1352 => to_slv(opcode_type, 16#11#),
      1353 => to_slv(opcode_type, 16#0F#),
      1354 => to_slv(opcode_type, 16#06#),
      1355 => to_slv(opcode_type, 16#0B#),
      1356 => to_slv(opcode_type, 16#56#),
      1357 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#08#),
      1377 => to_slv(opcode_type, 16#01#),
      1378 => to_slv(opcode_type, 16#03#),
      1379 => to_slv(opcode_type, 16#04#),
      1380 => to_slv(opcode_type, 16#9B#),
      1381 => to_slv(opcode_type, 16#03#),
      1382 => to_slv(opcode_type, 16#06#),
      1383 => to_slv(opcode_type, 16#08#),
      1384 => to_slv(opcode_type, 16#0A#),
      1385 => to_slv(opcode_type, 16#0E#),
      1386 => to_slv(opcode_type, 16#08#),
      1387 => to_slv(opcode_type, 16#11#),
      1388 => to_slv(opcode_type, 16#0E#),
      1389 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#07#),
      1409 => to_slv(opcode_type, 16#05#),
      1410 => to_slv(opcode_type, 16#09#),
      1411 => to_slv(opcode_type, 16#07#),
      1412 => to_slv(opcode_type, 16#10#),
      1413 => to_slv(opcode_type, 16#11#),
      1414 => to_slv(opcode_type, 16#01#),
      1415 => to_slv(opcode_type, 16#10#),
      1416 => to_slv(opcode_type, 16#03#),
      1417 => to_slv(opcode_type, 16#04#),
      1418 => to_slv(opcode_type, 16#06#),
      1419 => to_slv(opcode_type, 16#0B#),
      1420 => to_slv(opcode_type, 16#9A#),
      1421 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#04#),
      1441 => to_slv(opcode_type, 16#08#),
      1442 => to_slv(opcode_type, 16#01#),
      1443 => to_slv(opcode_type, 16#07#),
      1444 => to_slv(opcode_type, 16#11#),
      1445 => to_slv(opcode_type, 16#0C#),
      1446 => to_slv(opcode_type, 16#07#),
      1447 => to_slv(opcode_type, 16#07#),
      1448 => to_slv(opcode_type, 16#0D#),
      1449 => to_slv(opcode_type, 16#0F#),
      1450 => to_slv(opcode_type, 16#06#),
      1451 => to_slv(opcode_type, 16#0A#),
      1452 => to_slv(opcode_type, 16#0C#),
      1453 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#04#),
      1473 => to_slv(opcode_type, 16#07#),
      1474 => to_slv(opcode_type, 16#02#),
      1475 => to_slv(opcode_type, 16#09#),
      1476 => to_slv(opcode_type, 16#10#),
      1477 => to_slv(opcode_type, 16#0A#),
      1478 => to_slv(opcode_type, 16#06#),
      1479 => to_slv(opcode_type, 16#08#),
      1480 => to_slv(opcode_type, 16#0A#),
      1481 => to_slv(opcode_type, 16#0D#),
      1482 => to_slv(opcode_type, 16#08#),
      1483 => to_slv(opcode_type, 16#11#),
      1484 => to_slv(opcode_type, 16#0F#),
      1485 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#07#),
      1505 => to_slv(opcode_type, 16#05#),
      1506 => to_slv(opcode_type, 16#09#),
      1507 => to_slv(opcode_type, 16#04#),
      1508 => to_slv(opcode_type, 16#11#),
      1509 => to_slv(opcode_type, 16#04#),
      1510 => to_slv(opcode_type, 16#11#),
      1511 => to_slv(opcode_type, 16#06#),
      1512 => to_slv(opcode_type, 16#09#),
      1513 => to_slv(opcode_type, 16#04#),
      1514 => to_slv(opcode_type, 16#11#),
      1515 => to_slv(opcode_type, 16#0E#),
      1516 => to_slv(opcode_type, 16#0B#),
      1517 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#07#),
      1537 => to_slv(opcode_type, 16#03#),
      1538 => to_slv(opcode_type, 16#08#),
      1539 => to_slv(opcode_type, 16#03#),
      1540 => to_slv(opcode_type, 16#0A#),
      1541 => to_slv(opcode_type, 16#02#),
      1542 => to_slv(opcode_type, 16#0A#),
      1543 => to_slv(opcode_type, 16#01#),
      1544 => to_slv(opcode_type, 16#06#),
      1545 => to_slv(opcode_type, 16#02#),
      1546 => to_slv(opcode_type, 16#0F#),
      1547 => to_slv(opcode_type, 16#04#),
      1548 => to_slv(opcode_type, 16#0D#),
      1549 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#03#),
      1569 => to_slv(opcode_type, 16#09#),
      1570 => to_slv(opcode_type, 16#01#),
      1571 => to_slv(opcode_type, 16#09#),
      1572 => to_slv(opcode_type, 16#11#),
      1573 => to_slv(opcode_type, 16#10#),
      1574 => to_slv(opcode_type, 16#08#),
      1575 => to_slv(opcode_type, 16#07#),
      1576 => to_slv(opcode_type, 16#0F#),
      1577 => to_slv(opcode_type, 16#3A#),
      1578 => to_slv(opcode_type, 16#09#),
      1579 => to_slv(opcode_type, 16#0A#),
      1580 => to_slv(opcode_type, 16#0E#),
      1581 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#07#),
      1601 => to_slv(opcode_type, 16#09#),
      1602 => to_slv(opcode_type, 16#01#),
      1603 => to_slv(opcode_type, 16#09#),
      1604 => to_slv(opcode_type, 16#0D#),
      1605 => to_slv(opcode_type, 16#11#),
      1606 => to_slv(opcode_type, 16#03#),
      1607 => to_slv(opcode_type, 16#08#),
      1608 => to_slv(opcode_type, 16#0C#),
      1609 => to_slv(opcode_type, 16#63#),
      1610 => to_slv(opcode_type, 16#06#),
      1611 => to_slv(opcode_type, 16#0F#),
      1612 => to_slv(opcode_type, 16#0D#),
      1613 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#03#),
      1633 => to_slv(opcode_type, 16#07#),
      1634 => to_slv(opcode_type, 16#01#),
      1635 => to_slv(opcode_type, 16#06#),
      1636 => to_slv(opcode_type, 16#11#),
      1637 => to_slv(opcode_type, 16#11#),
      1638 => to_slv(opcode_type, 16#09#),
      1639 => to_slv(opcode_type, 16#06#),
      1640 => to_slv(opcode_type, 16#0C#),
      1641 => to_slv(opcode_type, 16#0F#),
      1642 => to_slv(opcode_type, 16#08#),
      1643 => to_slv(opcode_type, 16#0D#),
      1644 => to_slv(opcode_type, 16#0F#),
      1645 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#08#),
      1665 => to_slv(opcode_type, 16#03#),
      1666 => to_slv(opcode_type, 16#04#),
      1667 => to_slv(opcode_type, 16#01#),
      1668 => to_slv(opcode_type, 16#0A#),
      1669 => to_slv(opcode_type, 16#02#),
      1670 => to_slv(opcode_type, 16#08#),
      1671 => to_slv(opcode_type, 16#06#),
      1672 => to_slv(opcode_type, 16#0B#),
      1673 => to_slv(opcode_type, 16#11#),
      1674 => to_slv(opcode_type, 16#06#),
      1675 => to_slv(opcode_type, 16#0C#),
      1676 => to_slv(opcode_type, 16#0F#),
      1677 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#01#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#08#),
      1699 => to_slv(opcode_type, 16#08#),
      1700 => to_slv(opcode_type, 16#FA#),
      1701 => to_slv(opcode_type, 16#0E#),
      1702 => to_slv(opcode_type, 16#08#),
      1703 => to_slv(opcode_type, 16#0A#),
      1704 => to_slv(opcode_type, 16#10#),
      1705 => to_slv(opcode_type, 16#05#),
      1706 => to_slv(opcode_type, 16#08#),
      1707 => to_slv(opcode_type, 16#91#),
      1708 => to_slv(opcode_type, 16#0F#),
      1709 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#04#),
      1729 => to_slv(opcode_type, 16#06#),
      1730 => to_slv(opcode_type, 16#02#),
      1731 => to_slv(opcode_type, 16#06#),
      1732 => to_slv(opcode_type, 16#0A#),
      1733 => to_slv(opcode_type, 16#0A#),
      1734 => to_slv(opcode_type, 16#07#),
      1735 => to_slv(opcode_type, 16#06#),
      1736 => to_slv(opcode_type, 16#0F#),
      1737 => to_slv(opcode_type, 16#10#),
      1738 => to_slv(opcode_type, 16#08#),
      1739 => to_slv(opcode_type, 16#61#),
      1740 => to_slv(opcode_type, 16#56#),
      1741 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#07#),
      1761 => to_slv(opcode_type, 16#08#),
      1762 => to_slv(opcode_type, 16#08#),
      1763 => to_slv(opcode_type, 16#01#),
      1764 => to_slv(opcode_type, 16#0A#),
      1765 => to_slv(opcode_type, 16#07#),
      1766 => to_slv(opcode_type, 16#0E#),
      1767 => to_slv(opcode_type, 16#0C#),
      1768 => to_slv(opcode_type, 16#05#),
      1769 => to_slv(opcode_type, 16#04#),
      1770 => to_slv(opcode_type, 16#11#),
      1771 => to_slv(opcode_type, 16#02#),
      1772 => to_slv(opcode_type, 16#10#),
      1773 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#08#),
      1793 => to_slv(opcode_type, 16#09#),
      1794 => to_slv(opcode_type, 16#02#),
      1795 => to_slv(opcode_type, 16#03#),
      1796 => to_slv(opcode_type, 16#0C#),
      1797 => to_slv(opcode_type, 16#09#),
      1798 => to_slv(opcode_type, 16#03#),
      1799 => to_slv(opcode_type, 16#0D#),
      1800 => to_slv(opcode_type, 16#03#),
      1801 => to_slv(opcode_type, 16#0D#),
      1802 => to_slv(opcode_type, 16#04#),
      1803 => to_slv(opcode_type, 16#05#),
      1804 => to_slv(opcode_type, 16#B8#),
      1805 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#06#),
      1825 => to_slv(opcode_type, 16#03#),
      1826 => to_slv(opcode_type, 16#04#),
      1827 => to_slv(opcode_type, 16#08#),
      1828 => to_slv(opcode_type, 16#0F#),
      1829 => to_slv(opcode_type, 16#0C#),
      1830 => to_slv(opcode_type, 16#02#),
      1831 => to_slv(opcode_type, 16#09#),
      1832 => to_slv(opcode_type, 16#08#),
      1833 => to_slv(opcode_type, 16#0E#),
      1834 => to_slv(opcode_type, 16#10#),
      1835 => to_slv(opcode_type, 16#01#),
      1836 => to_slv(opcode_type, 16#0E#),
      1837 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#01#),
      1857 => to_slv(opcode_type, 16#06#),
      1858 => to_slv(opcode_type, 16#05#),
      1859 => to_slv(opcode_type, 16#07#),
      1860 => to_slv(opcode_type, 16#0B#),
      1861 => to_slv(opcode_type, 16#0F#),
      1862 => to_slv(opcode_type, 16#09#),
      1863 => to_slv(opcode_type, 16#06#),
      1864 => to_slv(opcode_type, 16#10#),
      1865 => to_slv(opcode_type, 16#0E#),
      1866 => to_slv(opcode_type, 16#08#),
      1867 => to_slv(opcode_type, 16#0F#),
      1868 => to_slv(opcode_type, 16#0A#),
      1869 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#05#),
      1889 => to_slv(opcode_type, 16#07#),
      1890 => to_slv(opcode_type, 16#02#),
      1891 => to_slv(opcode_type, 16#06#),
      1892 => to_slv(opcode_type, 16#0D#),
      1893 => to_slv(opcode_type, 16#0D#),
      1894 => to_slv(opcode_type, 16#07#),
      1895 => to_slv(opcode_type, 16#09#),
      1896 => to_slv(opcode_type, 16#0A#),
      1897 => to_slv(opcode_type, 16#0A#),
      1898 => to_slv(opcode_type, 16#06#),
      1899 => to_slv(opcode_type, 16#8E#),
      1900 => to_slv(opcode_type, 16#0A#),
      1901 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#08#),
      1921 => to_slv(opcode_type, 16#09#),
      1922 => to_slv(opcode_type, 16#08#),
      1923 => to_slv(opcode_type, 16#03#),
      1924 => to_slv(opcode_type, 16#0B#),
      1925 => to_slv(opcode_type, 16#09#),
      1926 => to_slv(opcode_type, 16#0C#),
      1927 => to_slv(opcode_type, 16#0B#),
      1928 => to_slv(opcode_type, 16#06#),
      1929 => to_slv(opcode_type, 16#03#),
      1930 => to_slv(opcode_type, 16#10#),
      1931 => to_slv(opcode_type, 16#59#),
      1932 => to_slv(opcode_type, 16#0A#),
      1933 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#09#),
      1953 => to_slv(opcode_type, 16#04#),
      1954 => to_slv(opcode_type, 16#03#),
      1955 => to_slv(opcode_type, 16#08#),
      1956 => to_slv(opcode_type, 16#0F#),
      1957 => to_slv(opcode_type, 16#0F#),
      1958 => to_slv(opcode_type, 16#03#),
      1959 => to_slv(opcode_type, 16#07#),
      1960 => to_slv(opcode_type, 16#05#),
      1961 => to_slv(opcode_type, 16#0D#),
      1962 => to_slv(opcode_type, 16#08#),
      1963 => to_slv(opcode_type, 16#0E#),
      1964 => to_slv(opcode_type, 16#0A#),
      1965 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#04#),
      1985 => to_slv(opcode_type, 16#09#),
      1986 => to_slv(opcode_type, 16#07#),
      1987 => to_slv(opcode_type, 16#05#),
      1988 => to_slv(opcode_type, 16#0C#),
      1989 => to_slv(opcode_type, 16#09#),
      1990 => to_slv(opcode_type, 16#11#),
      1991 => to_slv(opcode_type, 16#0D#),
      1992 => to_slv(opcode_type, 16#09#),
      1993 => to_slv(opcode_type, 16#02#),
      1994 => to_slv(opcode_type, 16#13#),
      1995 => to_slv(opcode_type, 16#03#),
      1996 => to_slv(opcode_type, 16#0F#),
      1997 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#02#),
      2017 => to_slv(opcode_type, 16#07#),
      2018 => to_slv(opcode_type, 16#03#),
      2019 => to_slv(opcode_type, 16#08#),
      2020 => to_slv(opcode_type, 16#14#),
      2021 => to_slv(opcode_type, 16#0A#),
      2022 => to_slv(opcode_type, 16#06#),
      2023 => to_slv(opcode_type, 16#06#),
      2024 => to_slv(opcode_type, 16#0E#),
      2025 => to_slv(opcode_type, 16#0B#),
      2026 => to_slv(opcode_type, 16#08#),
      2027 => to_slv(opcode_type, 16#0F#),
      2028 => to_slv(opcode_type, 16#24#),
      2029 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#03#),
      2049 => to_slv(opcode_type, 16#08#),
      2050 => to_slv(opcode_type, 16#08#),
      2051 => to_slv(opcode_type, 16#08#),
      2052 => to_slv(opcode_type, 16#CE#),
      2053 => to_slv(opcode_type, 16#0E#),
      2054 => to_slv(opcode_type, 16#07#),
      2055 => to_slv(opcode_type, 16#A1#),
      2056 => to_slv(opcode_type, 16#0D#),
      2057 => to_slv(opcode_type, 16#06#),
      2058 => to_slv(opcode_type, 16#04#),
      2059 => to_slv(opcode_type, 16#11#),
      2060 => to_slv(opcode_type, 16#0A#),
      2061 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#05#),
      2081 => to_slv(opcode_type, 16#09#),
      2082 => to_slv(opcode_type, 16#01#),
      2083 => to_slv(opcode_type, 16#07#),
      2084 => to_slv(opcode_type, 16#0B#),
      2085 => to_slv(opcode_type, 16#0C#),
      2086 => to_slv(opcode_type, 16#07#),
      2087 => to_slv(opcode_type, 16#09#),
      2088 => to_slv(opcode_type, 16#0D#),
      2089 => to_slv(opcode_type, 16#0F#),
      2090 => to_slv(opcode_type, 16#08#),
      2091 => to_slv(opcode_type, 16#11#),
      2092 => to_slv(opcode_type, 16#0E#),
      2093 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#02#),
      2113 => to_slv(opcode_type, 16#07#),
      2114 => to_slv(opcode_type, 16#05#),
      2115 => to_slv(opcode_type, 16#09#),
      2116 => to_slv(opcode_type, 16#0E#),
      2117 => to_slv(opcode_type, 16#0F#),
      2118 => to_slv(opcode_type, 16#08#),
      2119 => to_slv(opcode_type, 16#07#),
      2120 => to_slv(opcode_type, 16#0A#),
      2121 => to_slv(opcode_type, 16#10#),
      2122 => to_slv(opcode_type, 16#06#),
      2123 => to_slv(opcode_type, 16#11#),
      2124 => to_slv(opcode_type, 16#E2#),
      2125 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#05#),
      2145 => to_slv(opcode_type, 16#06#),
      2146 => to_slv(opcode_type, 16#04#),
      2147 => to_slv(opcode_type, 16#07#),
      2148 => to_slv(opcode_type, 16#78#),
      2149 => to_slv(opcode_type, 16#10#),
      2150 => to_slv(opcode_type, 16#08#),
      2151 => to_slv(opcode_type, 16#08#),
      2152 => to_slv(opcode_type, 16#24#),
      2153 => to_slv(opcode_type, 16#10#),
      2154 => to_slv(opcode_type, 16#06#),
      2155 => to_slv(opcode_type, 16#0B#),
      2156 => to_slv(opcode_type, 16#0D#),
      2157 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#02#),
      2177 => to_slv(opcode_type, 16#08#),
      2178 => to_slv(opcode_type, 16#07#),
      2179 => to_slv(opcode_type, 16#04#),
      2180 => to_slv(opcode_type, 16#0B#),
      2181 => to_slv(opcode_type, 16#09#),
      2182 => to_slv(opcode_type, 16#44#),
      2183 => to_slv(opcode_type, 16#10#),
      2184 => to_slv(opcode_type, 16#06#),
      2185 => to_slv(opcode_type, 16#04#),
      2186 => to_slv(opcode_type, 16#0C#),
      2187 => to_slv(opcode_type, 16#05#),
      2188 => to_slv(opcode_type, 16#11#),
      2189 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#01#),
      2209 => to_slv(opcode_type, 16#07#),
      2210 => to_slv(opcode_type, 16#03#),
      2211 => to_slv(opcode_type, 16#06#),
      2212 => to_slv(opcode_type, 16#0E#),
      2213 => to_slv(opcode_type, 16#10#),
      2214 => to_slv(opcode_type, 16#07#),
      2215 => to_slv(opcode_type, 16#06#),
      2216 => to_slv(opcode_type, 16#0A#),
      2217 => to_slv(opcode_type, 16#0B#),
      2218 => to_slv(opcode_type, 16#09#),
      2219 => to_slv(opcode_type, 16#DF#),
      2220 => to_slv(opcode_type, 16#58#),
      2221 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#05#),
      2241 => to_slv(opcode_type, 16#09#),
      2242 => to_slv(opcode_type, 16#06#),
      2243 => to_slv(opcode_type, 16#04#),
      2244 => to_slv(opcode_type, 16#0A#),
      2245 => to_slv(opcode_type, 16#08#),
      2246 => to_slv(opcode_type, 16#11#),
      2247 => to_slv(opcode_type, 16#89#),
      2248 => to_slv(opcode_type, 16#06#),
      2249 => to_slv(opcode_type, 16#06#),
      2250 => to_slv(opcode_type, 16#0C#),
      2251 => to_slv(opcode_type, 16#0F#),
      2252 => to_slv(opcode_type, 16#0B#),
      2253 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#09#),
      2273 => to_slv(opcode_type, 16#06#),
      2274 => to_slv(opcode_type, 16#05#),
      2275 => to_slv(opcode_type, 16#02#),
      2276 => to_slv(opcode_type, 16#0B#),
      2277 => to_slv(opcode_type, 16#09#),
      2278 => to_slv(opcode_type, 16#09#),
      2279 => to_slv(opcode_type, 16#0C#),
      2280 => to_slv(opcode_type, 16#0B#),
      2281 => to_slv(opcode_type, 16#02#),
      2282 => to_slv(opcode_type, 16#0C#),
      2283 => to_slv(opcode_type, 16#02#),
      2284 => to_slv(opcode_type, 16#0B#),
      2285 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#03#),
      2305 => to_slv(opcode_type, 16#07#),
      2306 => to_slv(opcode_type, 16#02#),
      2307 => to_slv(opcode_type, 16#08#),
      2308 => to_slv(opcode_type, 16#55#),
      2309 => to_slv(opcode_type, 16#10#),
      2310 => to_slv(opcode_type, 16#06#),
      2311 => to_slv(opcode_type, 16#06#),
      2312 => to_slv(opcode_type, 16#10#),
      2313 => to_slv(opcode_type, 16#0B#),
      2314 => to_slv(opcode_type, 16#07#),
      2315 => to_slv(opcode_type, 16#0A#),
      2316 => to_slv(opcode_type, 16#AF#),
      2317 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#07#),
      2337 => to_slv(opcode_type, 16#07#),
      2338 => to_slv(opcode_type, 16#02#),
      2339 => to_slv(opcode_type, 16#05#),
      2340 => to_slv(opcode_type, 16#0C#),
      2341 => to_slv(opcode_type, 16#06#),
      2342 => to_slv(opcode_type, 16#07#),
      2343 => to_slv(opcode_type, 16#11#),
      2344 => to_slv(opcode_type, 16#0F#),
      2345 => to_slv(opcode_type, 16#01#),
      2346 => to_slv(opcode_type, 16#0B#),
      2347 => to_slv(opcode_type, 16#01#),
      2348 => to_slv(opcode_type, 16#0A#),
      2349 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#04#),
      2369 => to_slv(opcode_type, 16#07#),
      2370 => to_slv(opcode_type, 16#09#),
      2371 => to_slv(opcode_type, 16#01#),
      2372 => to_slv(opcode_type, 16#0C#),
      2373 => to_slv(opcode_type, 16#06#),
      2374 => to_slv(opcode_type, 16#10#),
      2375 => to_slv(opcode_type, 16#0F#),
      2376 => to_slv(opcode_type, 16#07#),
      2377 => to_slv(opcode_type, 16#04#),
      2378 => to_slv(opcode_type, 16#0B#),
      2379 => to_slv(opcode_type, 16#05#),
      2380 => to_slv(opcode_type, 16#0F#),
      2381 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#07#),
      2401 => to_slv(opcode_type, 16#09#),
      2402 => to_slv(opcode_type, 16#05#),
      2403 => to_slv(opcode_type, 16#06#),
      2404 => to_slv(opcode_type, 16#0B#),
      2405 => to_slv(opcode_type, 16#11#),
      2406 => to_slv(opcode_type, 16#02#),
      2407 => to_slv(opcode_type, 16#06#),
      2408 => to_slv(opcode_type, 16#D9#),
      2409 => to_slv(opcode_type, 16#0C#),
      2410 => to_slv(opcode_type, 16#04#),
      2411 => to_slv(opcode_type, 16#03#),
      2412 => to_slv(opcode_type, 16#0E#),
      2413 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#08#),
      2433 => to_slv(opcode_type, 16#09#),
      2434 => to_slv(opcode_type, 16#06#),
      2435 => to_slv(opcode_type, 16#03#),
      2436 => to_slv(opcode_type, 16#0F#),
      2437 => to_slv(opcode_type, 16#06#),
      2438 => to_slv(opcode_type, 16#0F#),
      2439 => to_slv(opcode_type, 16#11#),
      2440 => to_slv(opcode_type, 16#09#),
      2441 => to_slv(opcode_type, 16#04#),
      2442 => to_slv(opcode_type, 16#11#),
      2443 => to_slv(opcode_type, 16#0C#),
      2444 => to_slv(opcode_type, 16#0B#),
      2445 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#03#),
      2465 => to_slv(opcode_type, 16#07#),
      2466 => to_slv(opcode_type, 16#03#),
      2467 => to_slv(opcode_type, 16#09#),
      2468 => to_slv(opcode_type, 16#0F#),
      2469 => to_slv(opcode_type, 16#12#),
      2470 => to_slv(opcode_type, 16#09#),
      2471 => to_slv(opcode_type, 16#09#),
      2472 => to_slv(opcode_type, 16#0E#),
      2473 => to_slv(opcode_type, 16#10#),
      2474 => to_slv(opcode_type, 16#07#),
      2475 => to_slv(opcode_type, 16#1B#),
      2476 => to_slv(opcode_type, 16#10#),
      2477 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#09#),
      2497 => to_slv(opcode_type, 16#03#),
      2498 => to_slv(opcode_type, 16#03#),
      2499 => to_slv(opcode_type, 16#09#),
      2500 => to_slv(opcode_type, 16#10#),
      2501 => to_slv(opcode_type, 16#0D#),
      2502 => to_slv(opcode_type, 16#01#),
      2503 => to_slv(opcode_type, 16#08#),
      2504 => to_slv(opcode_type, 16#06#),
      2505 => to_slv(opcode_type, 16#11#),
      2506 => to_slv(opcode_type, 16#0A#),
      2507 => to_slv(opcode_type, 16#04#),
      2508 => to_slv(opcode_type, 16#0C#),
      2509 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#02#),
      2529 => to_slv(opcode_type, 16#08#),
      2530 => to_slv(opcode_type, 16#04#),
      2531 => to_slv(opcode_type, 16#08#),
      2532 => to_slv(opcode_type, 16#0A#),
      2533 => to_slv(opcode_type, 16#11#),
      2534 => to_slv(opcode_type, 16#06#),
      2535 => to_slv(opcode_type, 16#08#),
      2536 => to_slv(opcode_type, 16#0A#),
      2537 => to_slv(opcode_type, 16#0D#),
      2538 => to_slv(opcode_type, 16#09#),
      2539 => to_slv(opcode_type, 16#11#),
      2540 => to_slv(opcode_type, 16#0E#),
      2541 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#08#),
      2561 => to_slv(opcode_type, 16#06#),
      2562 => to_slv(opcode_type, 16#01#),
      2563 => to_slv(opcode_type, 16#08#),
      2564 => to_slv(opcode_type, 16#0A#),
      2565 => to_slv(opcode_type, 16#10#),
      2566 => to_slv(opcode_type, 16#01#),
      2567 => to_slv(opcode_type, 16#03#),
      2568 => to_slv(opcode_type, 16#11#),
      2569 => to_slv(opcode_type, 16#04#),
      2570 => to_slv(opcode_type, 16#08#),
      2571 => to_slv(opcode_type, 16#FD#),
      2572 => to_slv(opcode_type, 16#0C#),
      2573 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#06#),
      2593 => to_slv(opcode_type, 16#02#),
      2594 => to_slv(opcode_type, 16#09#),
      2595 => to_slv(opcode_type, 16#02#),
      2596 => to_slv(opcode_type, 16#10#),
      2597 => to_slv(opcode_type, 16#02#),
      2598 => to_slv(opcode_type, 16#61#),
      2599 => to_slv(opcode_type, 16#09#),
      2600 => to_slv(opcode_type, 16#08#),
      2601 => to_slv(opcode_type, 16#03#),
      2602 => to_slv(opcode_type, 16#0F#),
      2603 => to_slv(opcode_type, 16#0A#),
      2604 => to_slv(opcode_type, 16#0C#),
      2605 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#03#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#09#),
      2627 => to_slv(opcode_type, 16#01#),
      2628 => to_slv(opcode_type, 16#0B#),
      2629 => to_slv(opcode_type, 16#08#),
      2630 => to_slv(opcode_type, 16#0A#),
      2631 => to_slv(opcode_type, 16#0A#),
      2632 => to_slv(opcode_type, 16#09#),
      2633 => to_slv(opcode_type, 16#07#),
      2634 => to_slv(opcode_type, 16#0E#),
      2635 => to_slv(opcode_type, 16#0A#),
      2636 => to_slv(opcode_type, 16#E3#),
      2637 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#04#),
      2657 => to_slv(opcode_type, 16#06#),
      2658 => to_slv(opcode_type, 16#05#),
      2659 => to_slv(opcode_type, 16#07#),
      2660 => to_slv(opcode_type, 16#0B#),
      2661 => to_slv(opcode_type, 16#0C#),
      2662 => to_slv(opcode_type, 16#06#),
      2663 => to_slv(opcode_type, 16#08#),
      2664 => to_slv(opcode_type, 16#0F#),
      2665 => to_slv(opcode_type, 16#0A#),
      2666 => to_slv(opcode_type, 16#09#),
      2667 => to_slv(opcode_type, 16#0F#),
      2668 => to_slv(opcode_type, 16#0B#),
      2669 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#08#),
      2689 => to_slv(opcode_type, 16#04#),
      2690 => to_slv(opcode_type, 16#03#),
      2691 => to_slv(opcode_type, 16#06#),
      2692 => to_slv(opcode_type, 16#10#),
      2693 => to_slv(opcode_type, 16#0E#),
      2694 => to_slv(opcode_type, 16#03#),
      2695 => to_slv(opcode_type, 16#09#),
      2696 => to_slv(opcode_type, 16#09#),
      2697 => to_slv(opcode_type, 16#0C#),
      2698 => to_slv(opcode_type, 16#10#),
      2699 => to_slv(opcode_type, 16#05#),
      2700 => to_slv(opcode_type, 16#0C#),
      2701 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#09#),
      2721 => to_slv(opcode_type, 16#04#),
      2722 => to_slv(opcode_type, 16#05#),
      2723 => to_slv(opcode_type, 16#08#),
      2724 => to_slv(opcode_type, 16#0D#),
      2725 => to_slv(opcode_type, 16#0C#),
      2726 => to_slv(opcode_type, 16#09#),
      2727 => to_slv(opcode_type, 16#02#),
      2728 => to_slv(opcode_type, 16#01#),
      2729 => to_slv(opcode_type, 16#0A#),
      2730 => to_slv(opcode_type, 16#05#),
      2731 => to_slv(opcode_type, 16#03#),
      2732 => to_slv(opcode_type, 16#0F#),
      2733 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#01#),
      2753 => to_slv(opcode_type, 16#08#),
      2754 => to_slv(opcode_type, 16#01#),
      2755 => to_slv(opcode_type, 16#09#),
      2756 => to_slv(opcode_type, 16#4F#),
      2757 => to_slv(opcode_type, 16#0A#),
      2758 => to_slv(opcode_type, 16#09#),
      2759 => to_slv(opcode_type, 16#08#),
      2760 => to_slv(opcode_type, 16#0A#),
      2761 => to_slv(opcode_type, 16#0C#),
      2762 => to_slv(opcode_type, 16#06#),
      2763 => to_slv(opcode_type, 16#10#),
      2764 => to_slv(opcode_type, 16#0A#),
      2765 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#05#),
      2785 => to_slv(opcode_type, 16#07#),
      2786 => to_slv(opcode_type, 16#02#),
      2787 => to_slv(opcode_type, 16#08#),
      2788 => to_slv(opcode_type, 16#0B#),
      2789 => to_slv(opcode_type, 16#10#),
      2790 => to_slv(opcode_type, 16#08#),
      2791 => to_slv(opcode_type, 16#08#),
      2792 => to_slv(opcode_type, 16#0A#),
      2793 => to_slv(opcode_type, 16#0B#),
      2794 => to_slv(opcode_type, 16#07#),
      2795 => to_slv(opcode_type, 16#0D#),
      2796 => to_slv(opcode_type, 16#0D#),
      2797 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#02#),
      2817 => to_slv(opcode_type, 16#08#),
      2818 => to_slv(opcode_type, 16#05#),
      2819 => to_slv(opcode_type, 16#08#),
      2820 => to_slv(opcode_type, 16#0A#),
      2821 => to_slv(opcode_type, 16#10#),
      2822 => to_slv(opcode_type, 16#08#),
      2823 => to_slv(opcode_type, 16#07#),
      2824 => to_slv(opcode_type, 16#0F#),
      2825 => to_slv(opcode_type, 16#0F#),
      2826 => to_slv(opcode_type, 16#09#),
      2827 => to_slv(opcode_type, 16#3A#),
      2828 => to_slv(opcode_type, 16#11#),
      2829 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#02#),
      2849 => to_slv(opcode_type, 16#09#),
      2850 => to_slv(opcode_type, 16#08#),
      2851 => to_slv(opcode_type, 16#07#),
      2852 => to_slv(opcode_type, 16#10#),
      2853 => to_slv(opcode_type, 16#0A#),
      2854 => to_slv(opcode_type, 16#04#),
      2855 => to_slv(opcode_type, 16#0E#),
      2856 => to_slv(opcode_type, 16#08#),
      2857 => to_slv(opcode_type, 16#06#),
      2858 => to_slv(opcode_type, 16#0E#),
      2859 => to_slv(opcode_type, 16#0A#),
      2860 => to_slv(opcode_type, 16#0F#),
      2861 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#02#),
      2881 => to_slv(opcode_type, 16#07#),
      2882 => to_slv(opcode_type, 16#02#),
      2883 => to_slv(opcode_type, 16#09#),
      2884 => to_slv(opcode_type, 16#0A#),
      2885 => to_slv(opcode_type, 16#0B#),
      2886 => to_slv(opcode_type, 16#06#),
      2887 => to_slv(opcode_type, 16#07#),
      2888 => to_slv(opcode_type, 16#11#),
      2889 => to_slv(opcode_type, 16#2B#),
      2890 => to_slv(opcode_type, 16#08#),
      2891 => to_slv(opcode_type, 16#0A#),
      2892 => to_slv(opcode_type, 16#0D#),
      2893 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#09#),
      2913 => to_slv(opcode_type, 16#09#),
      2914 => to_slv(opcode_type, 16#06#),
      2915 => to_slv(opcode_type, 16#07#),
      2916 => to_slv(opcode_type, 16#18#),
      2917 => to_slv(opcode_type, 16#0C#),
      2918 => to_slv(opcode_type, 16#09#),
      2919 => to_slv(opcode_type, 16#11#),
      2920 => to_slv(opcode_type, 16#0C#),
      2921 => to_slv(opcode_type, 16#09#),
      2922 => to_slv(opcode_type, 16#0B#),
      2923 => to_slv(opcode_type, 16#10#),
      2924 => to_slv(opcode_type, 16#11#),
      2925 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#09#),
      2945 => to_slv(opcode_type, 16#09#),
      2946 => to_slv(opcode_type, 16#08#),
      2947 => to_slv(opcode_type, 16#01#),
      2948 => to_slv(opcode_type, 16#0F#),
      2949 => to_slv(opcode_type, 16#08#),
      2950 => to_slv(opcode_type, 16#1D#),
      2951 => to_slv(opcode_type, 16#0E#),
      2952 => to_slv(opcode_type, 16#03#),
      2953 => to_slv(opcode_type, 16#02#),
      2954 => to_slv(opcode_type, 16#30#),
      2955 => to_slv(opcode_type, 16#05#),
      2956 => to_slv(opcode_type, 16#0C#),
      2957 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#04#),
      2977 => to_slv(opcode_type, 16#09#),
      2978 => to_slv(opcode_type, 16#05#),
      2979 => to_slv(opcode_type, 16#09#),
      2980 => to_slv(opcode_type, 16#0F#),
      2981 => to_slv(opcode_type, 16#11#),
      2982 => to_slv(opcode_type, 16#09#),
      2983 => to_slv(opcode_type, 16#09#),
      2984 => to_slv(opcode_type, 16#0D#),
      2985 => to_slv(opcode_type, 16#0E#),
      2986 => to_slv(opcode_type, 16#07#),
      2987 => to_slv(opcode_type, 16#0D#),
      2988 => to_slv(opcode_type, 16#0F#),
      2989 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#05#),
      3009 => to_slv(opcode_type, 16#09#),
      3010 => to_slv(opcode_type, 16#06#),
      3011 => to_slv(opcode_type, 16#09#),
      3012 => to_slv(opcode_type, 16#0C#),
      3013 => to_slv(opcode_type, 16#0D#),
      3014 => to_slv(opcode_type, 16#03#),
      3015 => to_slv(opcode_type, 16#0E#),
      3016 => to_slv(opcode_type, 16#09#),
      3017 => to_slv(opcode_type, 16#09#),
      3018 => to_slv(opcode_type, 16#0E#),
      3019 => to_slv(opcode_type, 16#0D#),
      3020 => to_slv(opcode_type, 16#0A#),
      3021 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#09#),
      3041 => to_slv(opcode_type, 16#06#),
      3042 => to_slv(opcode_type, 16#01#),
      3043 => to_slv(opcode_type, 16#02#),
      3044 => to_slv(opcode_type, 16#0B#),
      3045 => to_slv(opcode_type, 16#05#),
      3046 => to_slv(opcode_type, 16#09#),
      3047 => to_slv(opcode_type, 16#0D#),
      3048 => to_slv(opcode_type, 16#0C#),
      3049 => to_slv(opcode_type, 16#09#),
      3050 => to_slv(opcode_type, 16#01#),
      3051 => to_slv(opcode_type, 16#0D#),
      3052 => to_slv(opcode_type, 16#0B#),
      3053 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#01#),
      3073 => to_slv(opcode_type, 16#06#),
      3074 => to_slv(opcode_type, 16#07#),
      3075 => to_slv(opcode_type, 16#05#),
      3076 => to_slv(opcode_type, 16#10#),
      3077 => to_slv(opcode_type, 16#03#),
      3078 => to_slv(opcode_type, 16#0F#),
      3079 => to_slv(opcode_type, 16#08#),
      3080 => to_slv(opcode_type, 16#02#),
      3081 => to_slv(opcode_type, 16#0D#),
      3082 => to_slv(opcode_type, 16#07#),
      3083 => to_slv(opcode_type, 16#0A#),
      3084 => to_slv(opcode_type, 16#0E#),
      3085 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#02#),
      3105 => to_slv(opcode_type, 16#08#),
      3106 => to_slv(opcode_type, 16#02#),
      3107 => to_slv(opcode_type, 16#08#),
      3108 => to_slv(opcode_type, 16#11#),
      3109 => to_slv(opcode_type, 16#10#),
      3110 => to_slv(opcode_type, 16#07#),
      3111 => to_slv(opcode_type, 16#07#),
      3112 => to_slv(opcode_type, 16#0D#),
      3113 => to_slv(opcode_type, 16#10#),
      3114 => to_slv(opcode_type, 16#07#),
      3115 => to_slv(opcode_type, 16#0B#),
      3116 => to_slv(opcode_type, 16#0D#),
      3117 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#06#),
      3137 => to_slv(opcode_type, 16#08#),
      3138 => to_slv(opcode_type, 16#09#),
      3139 => to_slv(opcode_type, 16#01#),
      3140 => to_slv(opcode_type, 16#0D#),
      3141 => to_slv(opcode_type, 16#07#),
      3142 => to_slv(opcode_type, 16#10#),
      3143 => to_slv(opcode_type, 16#0D#),
      3144 => to_slv(opcode_type, 16#02#),
      3145 => to_slv(opcode_type, 16#03#),
      3146 => to_slv(opcode_type, 16#56#),
      3147 => to_slv(opcode_type, 16#05#),
      3148 => to_slv(opcode_type, 16#11#),
      3149 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#05#),
      3169 => to_slv(opcode_type, 16#08#),
      3170 => to_slv(opcode_type, 16#07#),
      3171 => to_slv(opcode_type, 16#07#),
      3172 => to_slv(opcode_type, 16#0F#),
      3173 => to_slv(opcode_type, 16#10#),
      3174 => to_slv(opcode_type, 16#05#),
      3175 => to_slv(opcode_type, 16#0A#),
      3176 => to_slv(opcode_type, 16#07#),
      3177 => to_slv(opcode_type, 16#09#),
      3178 => to_slv(opcode_type, 16#0C#),
      3179 => to_slv(opcode_type, 16#0F#),
      3180 => to_slv(opcode_type, 16#0A#),
      3181 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#03#),
      3201 => to_slv(opcode_type, 16#06#),
      3202 => to_slv(opcode_type, 16#09#),
      3203 => to_slv(opcode_type, 16#08#),
      3204 => to_slv(opcode_type, 16#0A#),
      3205 => to_slv(opcode_type, 16#0B#),
      3206 => to_slv(opcode_type, 16#03#),
      3207 => to_slv(opcode_type, 16#0B#),
      3208 => to_slv(opcode_type, 16#06#),
      3209 => to_slv(opcode_type, 16#05#),
      3210 => to_slv(opcode_type, 16#11#),
      3211 => to_slv(opcode_type, 16#01#),
      3212 => to_slv(opcode_type, 16#11#),
      3213 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#03#),
      3233 => to_slv(opcode_type, 16#08#),
      3234 => to_slv(opcode_type, 16#04#),
      3235 => to_slv(opcode_type, 16#08#),
      3236 => to_slv(opcode_type, 16#11#),
      3237 => to_slv(opcode_type, 16#0A#),
      3238 => to_slv(opcode_type, 16#06#),
      3239 => to_slv(opcode_type, 16#08#),
      3240 => to_slv(opcode_type, 16#0F#),
      3241 => to_slv(opcode_type, 16#11#),
      3242 => to_slv(opcode_type, 16#09#),
      3243 => to_slv(opcode_type, 16#0E#),
      3244 => to_slv(opcode_type, 16#0E#),
      3245 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#05#),
      3265 => to_slv(opcode_type, 16#08#),
      3266 => to_slv(opcode_type, 16#06#),
      3267 => to_slv(opcode_type, 16#04#),
      3268 => to_slv(opcode_type, 16#10#),
      3269 => to_slv(opcode_type, 16#01#),
      3270 => to_slv(opcode_type, 16#0A#),
      3271 => to_slv(opcode_type, 16#09#),
      3272 => to_slv(opcode_type, 16#06#),
      3273 => to_slv(opcode_type, 16#11#),
      3274 => to_slv(opcode_type, 16#0E#),
      3275 => to_slv(opcode_type, 16#05#),
      3276 => to_slv(opcode_type, 16#0A#),
      3277 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#02#),
      3297 => to_slv(opcode_type, 16#06#),
      3298 => to_slv(opcode_type, 16#02#),
      3299 => to_slv(opcode_type, 16#06#),
      3300 => to_slv(opcode_type, 16#0F#),
      3301 => to_slv(opcode_type, 16#10#),
      3302 => to_slv(opcode_type, 16#09#),
      3303 => to_slv(opcode_type, 16#06#),
      3304 => to_slv(opcode_type, 16#0F#),
      3305 => to_slv(opcode_type, 16#0E#),
      3306 => to_slv(opcode_type, 16#07#),
      3307 => to_slv(opcode_type, 16#10#),
      3308 => to_slv(opcode_type, 16#11#),
      3309 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#03#),
      3329 => to_slv(opcode_type, 16#07#),
      3330 => to_slv(opcode_type, 16#08#),
      3331 => to_slv(opcode_type, 16#04#),
      3332 => to_slv(opcode_type, 16#10#),
      3333 => to_slv(opcode_type, 16#06#),
      3334 => to_slv(opcode_type, 16#0B#),
      3335 => to_slv(opcode_type, 16#10#),
      3336 => to_slv(opcode_type, 16#06#),
      3337 => to_slv(opcode_type, 16#02#),
      3338 => to_slv(opcode_type, 16#0B#),
      3339 => to_slv(opcode_type, 16#04#),
      3340 => to_slv(opcode_type, 16#DC#),
      3341 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#09#),
      3361 => to_slv(opcode_type, 16#03#),
      3362 => to_slv(opcode_type, 16#01#),
      3363 => to_slv(opcode_type, 16#05#),
      3364 => to_slv(opcode_type, 16#0A#),
      3365 => to_slv(opcode_type, 16#07#),
      3366 => to_slv(opcode_type, 16#06#),
      3367 => to_slv(opcode_type, 16#01#),
      3368 => to_slv(opcode_type, 16#0F#),
      3369 => to_slv(opcode_type, 16#04#),
      3370 => to_slv(opcode_type, 16#0F#),
      3371 => to_slv(opcode_type, 16#01#),
      3372 => to_slv(opcode_type, 16#0B#),
      3373 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#06#),
      3393 => to_slv(opcode_type, 16#09#),
      3394 => to_slv(opcode_type, 16#09#),
      3395 => to_slv(opcode_type, 16#06#),
      3396 => to_slv(opcode_type, 16#0D#),
      3397 => to_slv(opcode_type, 16#0A#),
      3398 => to_slv(opcode_type, 16#04#),
      3399 => to_slv(opcode_type, 16#D6#),
      3400 => to_slv(opcode_type, 16#01#),
      3401 => to_slv(opcode_type, 16#01#),
      3402 => to_slv(opcode_type, 16#0E#),
      3403 => to_slv(opcode_type, 16#03#),
      3404 => to_slv(opcode_type, 16#0B#),
      3405 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#01#),
      3425 => to_slv(opcode_type, 16#07#),
      3426 => to_slv(opcode_type, 16#06#),
      3427 => to_slv(opcode_type, 16#04#),
      3428 => to_slv(opcode_type, 16#0F#),
      3429 => to_slv(opcode_type, 16#02#),
      3430 => to_slv(opcode_type, 16#0F#),
      3431 => to_slv(opcode_type, 16#06#),
      3432 => to_slv(opcode_type, 16#07#),
      3433 => to_slv(opcode_type, 16#0B#),
      3434 => to_slv(opcode_type, 16#0E#),
      3435 => to_slv(opcode_type, 16#05#),
      3436 => to_slv(opcode_type, 16#0B#),
      3437 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#03#),
      3457 => to_slv(opcode_type, 16#08#),
      3458 => to_slv(opcode_type, 16#02#),
      3459 => to_slv(opcode_type, 16#07#),
      3460 => to_slv(opcode_type, 16#11#),
      3461 => to_slv(opcode_type, 16#0B#),
      3462 => to_slv(opcode_type, 16#09#),
      3463 => to_slv(opcode_type, 16#09#),
      3464 => to_slv(opcode_type, 16#0B#),
      3465 => to_slv(opcode_type, 16#11#),
      3466 => to_slv(opcode_type, 16#09#),
      3467 => to_slv(opcode_type, 16#0E#),
      3468 => to_slv(opcode_type, 16#0F#),
      3469 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#04#),
      3489 => to_slv(opcode_type, 16#06#),
      3490 => to_slv(opcode_type, 16#05#),
      3491 => to_slv(opcode_type, 16#06#),
      3492 => to_slv(opcode_type, 16#0E#),
      3493 => to_slv(opcode_type, 16#63#),
      3494 => to_slv(opcode_type, 16#07#),
      3495 => to_slv(opcode_type, 16#07#),
      3496 => to_slv(opcode_type, 16#0B#),
      3497 => to_slv(opcode_type, 16#B6#),
      3498 => to_slv(opcode_type, 16#06#),
      3499 => to_slv(opcode_type, 16#0B#),
      3500 => to_slv(opcode_type, 16#0D#),
      3501 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#05#),
      3521 => to_slv(opcode_type, 16#06#),
      3522 => to_slv(opcode_type, 16#07#),
      3523 => to_slv(opcode_type, 16#08#),
      3524 => to_slv(opcode_type, 16#0E#),
      3525 => to_slv(opcode_type, 16#0C#),
      3526 => to_slv(opcode_type, 16#07#),
      3527 => to_slv(opcode_type, 16#0B#),
      3528 => to_slv(opcode_type, 16#FF#),
      3529 => to_slv(opcode_type, 16#07#),
      3530 => to_slv(opcode_type, 16#02#),
      3531 => to_slv(opcode_type, 16#11#),
      3532 => to_slv(opcode_type, 16#0B#),
      3533 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#07#),
      3553 => to_slv(opcode_type, 16#09#),
      3554 => to_slv(opcode_type, 16#02#),
      3555 => to_slv(opcode_type, 16#04#),
      3556 => to_slv(opcode_type, 16#0C#),
      3557 => to_slv(opcode_type, 16#02#),
      3558 => to_slv(opcode_type, 16#02#),
      3559 => to_slv(opcode_type, 16#0A#),
      3560 => to_slv(opcode_type, 16#09#),
      3561 => to_slv(opcode_type, 16#07#),
      3562 => to_slv(opcode_type, 16#0F#),
      3563 => to_slv(opcode_type, 16#0C#),
      3564 => to_slv(opcode_type, 16#0D#),
      3565 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#07#),
      3585 => to_slv(opcode_type, 16#06#),
      3586 => to_slv(opcode_type, 16#07#),
      3587 => to_slv(opcode_type, 16#05#),
      3588 => to_slv(opcode_type, 16#0C#),
      3589 => to_slv(opcode_type, 16#07#),
      3590 => to_slv(opcode_type, 16#0D#),
      3591 => to_slv(opcode_type, 16#0D#),
      3592 => to_slv(opcode_type, 16#02#),
      3593 => to_slv(opcode_type, 16#08#),
      3594 => to_slv(opcode_type, 16#10#),
      3595 => to_slv(opcode_type, 16#10#),
      3596 => to_slv(opcode_type, 16#0D#),
      3597 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#09#),
      3617 => to_slv(opcode_type, 16#05#),
      3618 => to_slv(opcode_type, 16#05#),
      3619 => to_slv(opcode_type, 16#06#),
      3620 => to_slv(opcode_type, 16#0D#),
      3621 => to_slv(opcode_type, 16#0B#),
      3622 => to_slv(opcode_type, 16#09#),
      3623 => to_slv(opcode_type, 16#08#),
      3624 => to_slv(opcode_type, 16#04#),
      3625 => to_slv(opcode_type, 16#0C#),
      3626 => to_slv(opcode_type, 16#05#),
      3627 => to_slv(opcode_type, 16#11#),
      3628 => to_slv(opcode_type, 16#A0#),
      3629 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#04#),
      3649 => to_slv(opcode_type, 16#09#),
      3650 => to_slv(opcode_type, 16#03#),
      3651 => to_slv(opcode_type, 16#07#),
      3652 => to_slv(opcode_type, 16#11#),
      3653 => to_slv(opcode_type, 16#0E#),
      3654 => to_slv(opcode_type, 16#07#),
      3655 => to_slv(opcode_type, 16#07#),
      3656 => to_slv(opcode_type, 16#0C#),
      3657 => to_slv(opcode_type, 16#0E#),
      3658 => to_slv(opcode_type, 16#06#),
      3659 => to_slv(opcode_type, 16#0A#),
      3660 => to_slv(opcode_type, 16#0A#),
      3661 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#08#),
      3681 => to_slv(opcode_type, 16#07#),
      3682 => to_slv(opcode_type, 16#08#),
      3683 => to_slv(opcode_type, 16#07#),
      3684 => to_slv(opcode_type, 16#0F#),
      3685 => to_slv(opcode_type, 16#0C#),
      3686 => to_slv(opcode_type, 16#02#),
      3687 => to_slv(opcode_type, 16#0C#),
      3688 => to_slv(opcode_type, 16#05#),
      3689 => to_slv(opcode_type, 16#04#),
      3690 => to_slv(opcode_type, 16#11#),
      3691 => to_slv(opcode_type, 16#05#),
      3692 => to_slv(opcode_type, 16#11#),
      3693 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#08#),
      3713 => to_slv(opcode_type, 16#09#),
      3714 => to_slv(opcode_type, 16#09#),
      3715 => to_slv(opcode_type, 16#08#),
      3716 => to_slv(opcode_type, 16#0B#),
      3717 => to_slv(opcode_type, 16#0F#),
      3718 => to_slv(opcode_type, 16#08#),
      3719 => to_slv(opcode_type, 16#0D#),
      3720 => to_slv(opcode_type, 16#0D#),
      3721 => to_slv(opcode_type, 16#02#),
      3722 => to_slv(opcode_type, 16#02#),
      3723 => to_slv(opcode_type, 16#0F#),
      3724 => to_slv(opcode_type, 16#11#),
      3725 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#08#),
      3745 => to_slv(opcode_type, 16#06#),
      3746 => to_slv(opcode_type, 16#04#),
      3747 => to_slv(opcode_type, 16#06#),
      3748 => to_slv(opcode_type, 16#0A#),
      3749 => to_slv(opcode_type, 16#0B#),
      3750 => to_slv(opcode_type, 16#04#),
      3751 => to_slv(opcode_type, 16#09#),
      3752 => to_slv(opcode_type, 16#2E#),
      3753 => to_slv(opcode_type, 16#A3#),
      3754 => to_slv(opcode_type, 16#06#),
      3755 => to_slv(opcode_type, 16#0A#),
      3756 => to_slv(opcode_type, 16#0B#),
      3757 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#01#),
      3777 => to_slv(opcode_type, 16#06#),
      3778 => to_slv(opcode_type, 16#01#),
      3779 => to_slv(opcode_type, 16#08#),
      3780 => to_slv(opcode_type, 16#0A#),
      3781 => to_slv(opcode_type, 16#0E#),
      3782 => to_slv(opcode_type, 16#07#),
      3783 => to_slv(opcode_type, 16#06#),
      3784 => to_slv(opcode_type, 16#11#),
      3785 => to_slv(opcode_type, 16#0E#),
      3786 => to_slv(opcode_type, 16#08#),
      3787 => to_slv(opcode_type, 16#10#),
      3788 => to_slv(opcode_type, 16#0E#),
      3789 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#06#),
      3809 => to_slv(opcode_type, 16#05#),
      3810 => to_slv(opcode_type, 16#01#),
      3811 => to_slv(opcode_type, 16#01#),
      3812 => to_slv(opcode_type, 16#0C#),
      3813 => to_slv(opcode_type, 16#08#),
      3814 => to_slv(opcode_type, 16#06#),
      3815 => to_slv(opcode_type, 16#04#),
      3816 => to_slv(opcode_type, 16#0E#),
      3817 => to_slv(opcode_type, 16#04#),
      3818 => to_slv(opcode_type, 16#0D#),
      3819 => to_slv(opcode_type, 16#03#),
      3820 => to_slv(opcode_type, 16#10#),
      3821 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#09#),
      3841 => to_slv(opcode_type, 16#08#),
      3842 => to_slv(opcode_type, 16#09#),
      3843 => to_slv(opcode_type, 16#02#),
      3844 => to_slv(opcode_type, 16#0A#),
      3845 => to_slv(opcode_type, 16#02#),
      3846 => to_slv(opcode_type, 16#3A#),
      3847 => to_slv(opcode_type, 16#01#),
      3848 => to_slv(opcode_type, 16#03#),
      3849 => to_slv(opcode_type, 16#0E#),
      3850 => to_slv(opcode_type, 16#02#),
      3851 => to_slv(opcode_type, 16#02#),
      3852 => to_slv(opcode_type, 16#0B#),
      3853 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#07#),
      3873 => to_slv(opcode_type, 16#05#),
      3874 => to_slv(opcode_type, 16#01#),
      3875 => to_slv(opcode_type, 16#05#),
      3876 => to_slv(opcode_type, 16#DF#),
      3877 => to_slv(opcode_type, 16#08#),
      3878 => to_slv(opcode_type, 16#09#),
      3879 => to_slv(opcode_type, 16#05#),
      3880 => to_slv(opcode_type, 16#11#),
      3881 => to_slv(opcode_type, 16#06#),
      3882 => to_slv(opcode_type, 16#0E#),
      3883 => to_slv(opcode_type, 16#0C#),
      3884 => to_slv(opcode_type, 16#0F#),
      3885 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#05#),
      3905 => to_slv(opcode_type, 16#09#),
      3906 => to_slv(opcode_type, 16#04#),
      3907 => to_slv(opcode_type, 16#07#),
      3908 => to_slv(opcode_type, 16#10#),
      3909 => to_slv(opcode_type, 16#0A#),
      3910 => to_slv(opcode_type, 16#06#),
      3911 => to_slv(opcode_type, 16#06#),
      3912 => to_slv(opcode_type, 16#11#),
      3913 => to_slv(opcode_type, 16#0C#),
      3914 => to_slv(opcode_type, 16#09#),
      3915 => to_slv(opcode_type, 16#0F#),
      3916 => to_slv(opcode_type, 16#0E#),
      3917 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#02#),
      3937 => to_slv(opcode_type, 16#09#),
      3938 => to_slv(opcode_type, 16#01#),
      3939 => to_slv(opcode_type, 16#06#),
      3940 => to_slv(opcode_type, 16#0E#),
      3941 => to_slv(opcode_type, 16#0E#),
      3942 => to_slv(opcode_type, 16#08#),
      3943 => to_slv(opcode_type, 16#08#),
      3944 => to_slv(opcode_type, 16#0D#),
      3945 => to_slv(opcode_type, 16#0D#),
      3946 => to_slv(opcode_type, 16#09#),
      3947 => to_slv(opcode_type, 16#3B#),
      3948 => to_slv(opcode_type, 16#0B#),
      3949 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#05#),
      3969 => to_slv(opcode_type, 16#06#),
      3970 => to_slv(opcode_type, 16#07#),
      3971 => to_slv(opcode_type, 16#02#),
      3972 => to_slv(opcode_type, 16#11#),
      3973 => to_slv(opcode_type, 16#05#),
      3974 => to_slv(opcode_type, 16#11#),
      3975 => to_slv(opcode_type, 16#06#),
      3976 => to_slv(opcode_type, 16#02#),
      3977 => to_slv(opcode_type, 16#11#),
      3978 => to_slv(opcode_type, 16#07#),
      3979 => to_slv(opcode_type, 16#11#),
      3980 => to_slv(opcode_type, 16#11#),
      3981 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#08#),
      4001 => to_slv(opcode_type, 16#09#),
      4002 => to_slv(opcode_type, 16#04#),
      4003 => to_slv(opcode_type, 16#02#),
      4004 => to_slv(opcode_type, 16#0B#),
      4005 => to_slv(opcode_type, 16#04#),
      4006 => to_slv(opcode_type, 16#09#),
      4007 => to_slv(opcode_type, 16#B4#),
      4008 => to_slv(opcode_type, 16#0E#),
      4009 => to_slv(opcode_type, 16#08#),
      4010 => to_slv(opcode_type, 16#02#),
      4011 => to_slv(opcode_type, 16#10#),
      4012 => to_slv(opcode_type, 16#0D#),
      4013 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#07#),
      4033 => to_slv(opcode_type, 16#07#),
      4034 => to_slv(opcode_type, 16#09#),
      4035 => to_slv(opcode_type, 16#06#),
      4036 => to_slv(opcode_type, 16#0C#),
      4037 => to_slv(opcode_type, 16#0C#),
      4038 => to_slv(opcode_type, 16#06#),
      4039 => to_slv(opcode_type, 16#0A#),
      4040 => to_slv(opcode_type, 16#0E#),
      4041 => to_slv(opcode_type, 16#09#),
      4042 => to_slv(opcode_type, 16#10#),
      4043 => to_slv(opcode_type, 16#10#),
      4044 => to_slv(opcode_type, 16#0B#),
      4045 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#05#),
      4066 => to_slv(opcode_type, 16#09#),
      4067 => to_slv(opcode_type, 16#05#),
      4068 => to_slv(opcode_type, 16#0E#),
      4069 => to_slv(opcode_type, 16#05#),
      4070 => to_slv(opcode_type, 16#49#),
      4071 => to_slv(opcode_type, 16#07#),
      4072 => to_slv(opcode_type, 16#08#),
      4073 => to_slv(opcode_type, 16#04#),
      4074 => to_slv(opcode_type, 16#0F#),
      4075 => to_slv(opcode_type, 16#0C#),
      4076 => to_slv(opcode_type, 16#0F#),
      4077 to 4095 => (others => '0')
  ),

    -- Bin `14`...
    13 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#03#),
      1 => to_slv(opcode_type, 16#08#),
      2 => to_slv(opcode_type, 16#06#),
      3 => to_slv(opcode_type, 16#01#),
      4 => to_slv(opcode_type, 16#10#),
      5 => to_slv(opcode_type, 16#06#),
      6 => to_slv(opcode_type, 16#0F#),
      7 => to_slv(opcode_type, 16#D6#),
      8 => to_slv(opcode_type, 16#08#),
      9 => to_slv(opcode_type, 16#03#),
      10 => to_slv(opcode_type, 16#11#),
      11 => to_slv(opcode_type, 16#09#),
      12 => to_slv(opcode_type, 16#0C#),
      13 => to_slv(opcode_type, 16#0E#),
      14 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#09#),
      33 => to_slv(opcode_type, 16#01#),
      34 => to_slv(opcode_type, 16#05#),
      35 => to_slv(opcode_type, 16#09#),
      36 => to_slv(opcode_type, 16#0E#),
      37 => to_slv(opcode_type, 16#0C#),
      38 => to_slv(opcode_type, 16#09#),
      39 => to_slv(opcode_type, 16#04#),
      40 => to_slv(opcode_type, 16#07#),
      41 => to_slv(opcode_type, 16#0F#),
      42 => to_slv(opcode_type, 16#0F#),
      43 => to_slv(opcode_type, 16#07#),
      44 => to_slv(opcode_type, 16#0D#),
      45 => to_slv(opcode_type, 16#0C#),
      46 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#02#),
      65 => to_slv(opcode_type, 16#06#),
      66 => to_slv(opcode_type, 16#06#),
      67 => to_slv(opcode_type, 16#03#),
      68 => to_slv(opcode_type, 16#10#),
      69 => to_slv(opcode_type, 16#01#),
      70 => to_slv(opcode_type, 16#11#),
      71 => to_slv(opcode_type, 16#08#),
      72 => to_slv(opcode_type, 16#06#),
      73 => to_slv(opcode_type, 16#0E#),
      74 => to_slv(opcode_type, 16#0D#),
      75 => to_slv(opcode_type, 16#07#),
      76 => to_slv(opcode_type, 16#0D#),
      77 => to_slv(opcode_type, 16#10#),
      78 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#03#),
      97 => to_slv(opcode_type, 16#07#),
      98 => to_slv(opcode_type, 16#06#),
      99 => to_slv(opcode_type, 16#06#),
      100 => to_slv(opcode_type, 16#10#),
      101 => to_slv(opcode_type, 16#0B#),
      102 => to_slv(opcode_type, 16#07#),
      103 => to_slv(opcode_type, 16#0B#),
      104 => to_slv(opcode_type, 16#0A#),
      105 => to_slv(opcode_type, 16#07#),
      106 => to_slv(opcode_type, 16#04#),
      107 => to_slv(opcode_type, 16#0B#),
      108 => to_slv(opcode_type, 16#02#),
      109 => to_slv(opcode_type, 16#0A#),
      110 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#05#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#09#),
      131 => to_slv(opcode_type, 16#05#),
      132 => to_slv(opcode_type, 16#0A#),
      133 => to_slv(opcode_type, 16#05#),
      134 => to_slv(opcode_type, 16#11#),
      135 => to_slv(opcode_type, 16#08#),
      136 => to_slv(opcode_type, 16#07#),
      137 => to_slv(opcode_type, 16#0A#),
      138 => to_slv(opcode_type, 16#3A#),
      139 => to_slv(opcode_type, 16#08#),
      140 => to_slv(opcode_type, 16#0B#),
      141 => to_slv(opcode_type, 16#11#),
      142 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#08#),
      161 => to_slv(opcode_type, 16#05#),
      162 => to_slv(opcode_type, 16#01#),
      163 => to_slv(opcode_type, 16#08#),
      164 => to_slv(opcode_type, 16#8B#),
      165 => to_slv(opcode_type, 16#0E#),
      166 => to_slv(opcode_type, 16#03#),
      167 => to_slv(opcode_type, 16#07#),
      168 => to_slv(opcode_type, 16#07#),
      169 => to_slv(opcode_type, 16#0E#),
      170 => to_slv(opcode_type, 16#0D#),
      171 => to_slv(opcode_type, 16#08#),
      172 => to_slv(opcode_type, 16#10#),
      173 => to_slv(opcode_type, 16#10#),
      174 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#03#),
      193 => to_slv(opcode_type, 16#08#),
      194 => to_slv(opcode_type, 16#07#),
      195 => to_slv(opcode_type, 16#04#),
      196 => to_slv(opcode_type, 16#11#),
      197 => to_slv(opcode_type, 16#03#),
      198 => to_slv(opcode_type, 16#0D#),
      199 => to_slv(opcode_type, 16#07#),
      200 => to_slv(opcode_type, 16#07#),
      201 => to_slv(opcode_type, 16#5A#),
      202 => to_slv(opcode_type, 16#0E#),
      203 => to_slv(opcode_type, 16#09#),
      204 => to_slv(opcode_type, 16#C8#),
      205 => to_slv(opcode_type, 16#11#),
      206 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#09#),
      225 => to_slv(opcode_type, 16#07#),
      226 => to_slv(opcode_type, 16#08#),
      227 => to_slv(opcode_type, 16#08#),
      228 => to_slv(opcode_type, 16#CF#),
      229 => to_slv(opcode_type, 16#0B#),
      230 => to_slv(opcode_type, 16#08#),
      231 => to_slv(opcode_type, 16#0E#),
      232 => to_slv(opcode_type, 16#0D#),
      233 => to_slv(opcode_type, 16#04#),
      234 => to_slv(opcode_type, 16#05#),
      235 => to_slv(opcode_type, 16#0D#),
      236 => to_slv(opcode_type, 16#04#),
      237 => to_slv(opcode_type, 16#0E#),
      238 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#07#),
      257 => to_slv(opcode_type, 16#01#),
      258 => to_slv(opcode_type, 16#02#),
      259 => to_slv(opcode_type, 16#08#),
      260 => to_slv(opcode_type, 16#83#),
      261 => to_slv(opcode_type, 16#0F#),
      262 => to_slv(opcode_type, 16#09#),
      263 => to_slv(opcode_type, 16#03#),
      264 => to_slv(opcode_type, 16#04#),
      265 => to_slv(opcode_type, 16#10#),
      266 => to_slv(opcode_type, 16#03#),
      267 => to_slv(opcode_type, 16#09#),
      268 => to_slv(opcode_type, 16#0A#),
      269 => to_slv(opcode_type, 16#11#),
      270 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#09#),
      289 => to_slv(opcode_type, 16#03#),
      290 => to_slv(opcode_type, 16#02#),
      291 => to_slv(opcode_type, 16#04#),
      292 => to_slv(opcode_type, 16#0C#),
      293 => to_slv(opcode_type, 16#06#),
      294 => to_slv(opcode_type, 16#05#),
      295 => to_slv(opcode_type, 16#08#),
      296 => to_slv(opcode_type, 16#10#),
      297 => to_slv(opcode_type, 16#0D#),
      298 => to_slv(opcode_type, 16#05#),
      299 => to_slv(opcode_type, 16#07#),
      300 => to_slv(opcode_type, 16#10#),
      301 => to_slv(opcode_type, 16#0E#),
      302 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#08#),
      321 => to_slv(opcode_type, 16#09#),
      322 => to_slv(opcode_type, 16#01#),
      323 => to_slv(opcode_type, 16#09#),
      324 => to_slv(opcode_type, 16#0B#),
      325 => to_slv(opcode_type, 16#11#),
      326 => to_slv(opcode_type, 16#05#),
      327 => to_slv(opcode_type, 16#03#),
      328 => to_slv(opcode_type, 16#10#),
      329 => to_slv(opcode_type, 16#09#),
      330 => to_slv(opcode_type, 16#09#),
      331 => to_slv(opcode_type, 16#3A#),
      332 => to_slv(opcode_type, 16#8C#),
      333 => to_slv(opcode_type, 16#0E#),
      334 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#02#),
      353 => to_slv(opcode_type, 16#07#),
      354 => to_slv(opcode_type, 16#08#),
      355 => to_slv(opcode_type, 16#04#),
      356 => to_slv(opcode_type, 16#0E#),
      357 => to_slv(opcode_type, 16#06#),
      358 => to_slv(opcode_type, 16#11#),
      359 => to_slv(opcode_type, 16#3F#),
      360 => to_slv(opcode_type, 16#06#),
      361 => to_slv(opcode_type, 16#02#),
      362 => to_slv(opcode_type, 16#B9#),
      363 => to_slv(opcode_type, 16#09#),
      364 => to_slv(opcode_type, 16#10#),
      365 => to_slv(opcode_type, 16#0C#),
      366 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#04#),
      385 => to_slv(opcode_type, 16#08#),
      386 => to_slv(opcode_type, 16#06#),
      387 => to_slv(opcode_type, 16#04#),
      388 => to_slv(opcode_type, 16#0A#),
      389 => to_slv(opcode_type, 16#02#),
      390 => to_slv(opcode_type, 16#0C#),
      391 => to_slv(opcode_type, 16#06#),
      392 => to_slv(opcode_type, 16#07#),
      393 => to_slv(opcode_type, 16#0A#),
      394 => to_slv(opcode_type, 16#0C#),
      395 => to_slv(opcode_type, 16#06#),
      396 => to_slv(opcode_type, 16#10#),
      397 => to_slv(opcode_type, 16#10#),
      398 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#07#),
      417 => to_slv(opcode_type, 16#01#),
      418 => to_slv(opcode_type, 16#04#),
      419 => to_slv(opcode_type, 16#09#),
      420 => to_slv(opcode_type, 16#F9#),
      421 => to_slv(opcode_type, 16#10#),
      422 => to_slv(opcode_type, 16#02#),
      423 => to_slv(opcode_type, 16#08#),
      424 => to_slv(opcode_type, 16#06#),
      425 => to_slv(opcode_type, 16#0F#),
      426 => to_slv(opcode_type, 16#0B#),
      427 => to_slv(opcode_type, 16#06#),
      428 => to_slv(opcode_type, 16#0B#),
      429 => to_slv(opcode_type, 16#0A#),
      430 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#07#),
      449 => to_slv(opcode_type, 16#02#),
      450 => to_slv(opcode_type, 16#09#),
      451 => to_slv(opcode_type, 16#08#),
      452 => to_slv(opcode_type, 16#0C#),
      453 => to_slv(opcode_type, 16#0B#),
      454 => to_slv(opcode_type, 16#02#),
      455 => to_slv(opcode_type, 16#6A#),
      456 => to_slv(opcode_type, 16#03#),
      457 => to_slv(opcode_type, 16#08#),
      458 => to_slv(opcode_type, 16#03#),
      459 => to_slv(opcode_type, 16#0C#),
      460 => to_slv(opcode_type, 16#03#),
      461 => to_slv(opcode_type, 16#0F#),
      462 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#02#),
      481 => to_slv(opcode_type, 16#08#),
      482 => to_slv(opcode_type, 16#06#),
      483 => to_slv(opcode_type, 16#08#),
      484 => to_slv(opcode_type, 16#0F#),
      485 => to_slv(opcode_type, 16#15#),
      486 => to_slv(opcode_type, 16#05#),
      487 => to_slv(opcode_type, 16#0E#),
      488 => to_slv(opcode_type, 16#07#),
      489 => to_slv(opcode_type, 16#09#),
      490 => to_slv(opcode_type, 16#0C#),
      491 => to_slv(opcode_type, 16#0C#),
      492 => to_slv(opcode_type, 16#04#),
      493 => to_slv(opcode_type, 16#0C#),
      494 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#02#),
      513 => to_slv(opcode_type, 16#08#),
      514 => to_slv(opcode_type, 16#07#),
      515 => to_slv(opcode_type, 16#02#),
      516 => to_slv(opcode_type, 16#0B#),
      517 => to_slv(opcode_type, 16#02#),
      518 => to_slv(opcode_type, 16#0A#),
      519 => to_slv(opcode_type, 16#09#),
      520 => to_slv(opcode_type, 16#09#),
      521 => to_slv(opcode_type, 16#11#),
      522 => to_slv(opcode_type, 16#0C#),
      523 => to_slv(opcode_type, 16#09#),
      524 => to_slv(opcode_type, 16#0E#),
      525 => to_slv(opcode_type, 16#11#),
      526 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#01#),
      545 => to_slv(opcode_type, 16#09#),
      546 => to_slv(opcode_type, 16#08#),
      547 => to_slv(opcode_type, 16#02#),
      548 => to_slv(opcode_type, 16#0F#),
      549 => to_slv(opcode_type, 16#09#),
      550 => to_slv(opcode_type, 16#10#),
      551 => to_slv(opcode_type, 16#0D#),
      552 => to_slv(opcode_type, 16#07#),
      553 => to_slv(opcode_type, 16#05#),
      554 => to_slv(opcode_type, 16#0B#),
      555 => to_slv(opcode_type, 16#08#),
      556 => to_slv(opcode_type, 16#0D#),
      557 => to_slv(opcode_type, 16#33#),
      558 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#06#),
      577 => to_slv(opcode_type, 16#03#),
      578 => to_slv(opcode_type, 16#02#),
      579 => to_slv(opcode_type, 16#02#),
      580 => to_slv(opcode_type, 16#0A#),
      581 => to_slv(opcode_type, 16#06#),
      582 => to_slv(opcode_type, 16#02#),
      583 => to_slv(opcode_type, 16#06#),
      584 => to_slv(opcode_type, 16#0C#),
      585 => to_slv(opcode_type, 16#0A#),
      586 => to_slv(opcode_type, 16#08#),
      587 => to_slv(opcode_type, 16#01#),
      588 => to_slv(opcode_type, 16#78#),
      589 => to_slv(opcode_type, 16#0E#),
      590 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#04#),
      609 => to_slv(opcode_type, 16#06#),
      610 => to_slv(opcode_type, 16#07#),
      611 => to_slv(opcode_type, 16#04#),
      612 => to_slv(opcode_type, 16#0B#),
      613 => to_slv(opcode_type, 16#04#),
      614 => to_slv(opcode_type, 16#0D#),
      615 => to_slv(opcode_type, 16#07#),
      616 => to_slv(opcode_type, 16#08#),
      617 => to_slv(opcode_type, 16#0F#),
      618 => to_slv(opcode_type, 16#0B#),
      619 => to_slv(opcode_type, 16#07#),
      620 => to_slv(opcode_type, 16#0A#),
      621 => to_slv(opcode_type, 16#0C#),
      622 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#04#),
      641 => to_slv(opcode_type, 16#09#),
      642 => to_slv(opcode_type, 16#08#),
      643 => to_slv(opcode_type, 16#03#),
      644 => to_slv(opcode_type, 16#11#),
      645 => to_slv(opcode_type, 16#07#),
      646 => to_slv(opcode_type, 16#0E#),
      647 => to_slv(opcode_type, 16#0B#),
      648 => to_slv(opcode_type, 16#09#),
      649 => to_slv(opcode_type, 16#05#),
      650 => to_slv(opcode_type, 16#0C#),
      651 => to_slv(opcode_type, 16#07#),
      652 => to_slv(opcode_type, 16#0A#),
      653 => to_slv(opcode_type, 16#0E#),
      654 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#09#),
      673 => to_slv(opcode_type, 16#01#),
      674 => to_slv(opcode_type, 16#06#),
      675 => to_slv(opcode_type, 16#06#),
      676 => to_slv(opcode_type, 16#53#),
      677 => to_slv(opcode_type, 16#0F#),
      678 => to_slv(opcode_type, 16#05#),
      679 => to_slv(opcode_type, 16#0F#),
      680 => to_slv(opcode_type, 16#09#),
      681 => to_slv(opcode_type, 16#05#),
      682 => to_slv(opcode_type, 16#07#),
      683 => to_slv(opcode_type, 16#11#),
      684 => to_slv(opcode_type, 16#87#),
      685 => to_slv(opcode_type, 16#79#),
      686 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#09#),
      705 => to_slv(opcode_type, 16#07#),
      706 => to_slv(opcode_type, 16#04#),
      707 => to_slv(opcode_type, 16#07#),
      708 => to_slv(opcode_type, 16#0D#),
      709 => to_slv(opcode_type, 16#0C#),
      710 => to_slv(opcode_type, 16#03#),
      711 => to_slv(opcode_type, 16#08#),
      712 => to_slv(opcode_type, 16#0D#),
      713 => to_slv(opcode_type, 16#11#),
      714 => to_slv(opcode_type, 16#02#),
      715 => to_slv(opcode_type, 16#03#),
      716 => to_slv(opcode_type, 16#03#),
      717 => to_slv(opcode_type, 16#0D#),
      718 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#06#),
      737 => to_slv(opcode_type, 16#06#),
      738 => to_slv(opcode_type, 16#09#),
      739 => to_slv(opcode_type, 16#01#),
      740 => to_slv(opcode_type, 16#10#),
      741 => to_slv(opcode_type, 16#04#),
      742 => to_slv(opcode_type, 16#0E#),
      743 => to_slv(opcode_type, 16#04#),
      744 => to_slv(opcode_type, 16#08#),
      745 => to_slv(opcode_type, 16#0E#),
      746 => to_slv(opcode_type, 16#11#),
      747 => to_slv(opcode_type, 16#03#),
      748 => to_slv(opcode_type, 16#04#),
      749 => to_slv(opcode_type, 16#11#),
      750 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#05#),
      769 => to_slv(opcode_type, 16#08#),
      770 => to_slv(opcode_type, 16#06#),
      771 => to_slv(opcode_type, 16#04#),
      772 => to_slv(opcode_type, 16#0B#),
      773 => to_slv(opcode_type, 16#05#),
      774 => to_slv(opcode_type, 16#47#),
      775 => to_slv(opcode_type, 16#09#),
      776 => to_slv(opcode_type, 16#06#),
      777 => to_slv(opcode_type, 16#0D#),
      778 => to_slv(opcode_type, 16#0B#),
      779 => to_slv(opcode_type, 16#09#),
      780 => to_slv(opcode_type, 16#10#),
      781 => to_slv(opcode_type, 16#0C#),
      782 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#09#),
      801 => to_slv(opcode_type, 16#04#),
      802 => to_slv(opcode_type, 16#08#),
      803 => to_slv(opcode_type, 16#03#),
      804 => to_slv(opcode_type, 16#0A#),
      805 => to_slv(opcode_type, 16#01#),
      806 => to_slv(opcode_type, 16#0A#),
      807 => to_slv(opcode_type, 16#09#),
      808 => to_slv(opcode_type, 16#01#),
      809 => to_slv(opcode_type, 16#09#),
      810 => to_slv(opcode_type, 16#0D#),
      811 => to_slv(opcode_type, 16#0E#),
      812 => to_slv(opcode_type, 16#03#),
      813 => to_slv(opcode_type, 16#0B#),
      814 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#06#),
      833 => to_slv(opcode_type, 16#03#),
      834 => to_slv(opcode_type, 16#01#),
      835 => to_slv(opcode_type, 16#03#),
      836 => to_slv(opcode_type, 16#0C#),
      837 => to_slv(opcode_type, 16#07#),
      838 => to_slv(opcode_type, 16#03#),
      839 => to_slv(opcode_type, 16#01#),
      840 => to_slv(opcode_type, 16#0F#),
      841 => to_slv(opcode_type, 16#08#),
      842 => to_slv(opcode_type, 16#01#),
      843 => to_slv(opcode_type, 16#0B#),
      844 => to_slv(opcode_type, 16#01#),
      845 => to_slv(opcode_type, 16#11#),
      846 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#01#),
      865 => to_slv(opcode_type, 16#06#),
      866 => to_slv(opcode_type, 16#06#),
      867 => to_slv(opcode_type, 16#04#),
      868 => to_slv(opcode_type, 16#0D#),
      869 => to_slv(opcode_type, 16#05#),
      870 => to_slv(opcode_type, 16#0B#),
      871 => to_slv(opcode_type, 16#09#),
      872 => to_slv(opcode_type, 16#06#),
      873 => to_slv(opcode_type, 16#10#),
      874 => to_slv(opcode_type, 16#0D#),
      875 => to_slv(opcode_type, 16#06#),
      876 => to_slv(opcode_type, 16#11#),
      877 => to_slv(opcode_type, 16#0E#),
      878 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#08#),
      897 => to_slv(opcode_type, 16#05#),
      898 => to_slv(opcode_type, 16#01#),
      899 => to_slv(opcode_type, 16#05#),
      900 => to_slv(opcode_type, 16#0D#),
      901 => to_slv(opcode_type, 16#06#),
      902 => to_slv(opcode_type, 16#02#),
      903 => to_slv(opcode_type, 16#04#),
      904 => to_slv(opcode_type, 16#0B#),
      905 => to_slv(opcode_type, 16#07#),
      906 => to_slv(opcode_type, 16#02#),
      907 => to_slv(opcode_type, 16#0A#),
      908 => to_slv(opcode_type, 16#03#),
      909 => to_slv(opcode_type, 16#0B#),
      910 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#08#),
      929 => to_slv(opcode_type, 16#01#),
      930 => to_slv(opcode_type, 16#08#),
      931 => to_slv(opcode_type, 16#01#),
      932 => to_slv(opcode_type, 16#0E#),
      933 => to_slv(opcode_type, 16#09#),
      934 => to_slv(opcode_type, 16#11#),
      935 => to_slv(opcode_type, 16#10#),
      936 => to_slv(opcode_type, 16#08#),
      937 => to_slv(opcode_type, 16#05#),
      938 => to_slv(opcode_type, 16#03#),
      939 => to_slv(opcode_type, 16#0F#),
      940 => to_slv(opcode_type, 16#01#),
      941 => to_slv(opcode_type, 16#9B#),
      942 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#03#),
      961 => to_slv(opcode_type, 16#06#),
      962 => to_slv(opcode_type, 16#08#),
      963 => to_slv(opcode_type, 16#05#),
      964 => to_slv(opcode_type, 16#0C#),
      965 => to_slv(opcode_type, 16#02#),
      966 => to_slv(opcode_type, 16#10#),
      967 => to_slv(opcode_type, 16#07#),
      968 => to_slv(opcode_type, 16#07#),
      969 => to_slv(opcode_type, 16#0C#),
      970 => to_slv(opcode_type, 16#10#),
      971 => to_slv(opcode_type, 16#06#),
      972 => to_slv(opcode_type, 16#0A#),
      973 => to_slv(opcode_type, 16#11#),
      974 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#01#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#06#),
      995 => to_slv(opcode_type, 16#08#),
      996 => to_slv(opcode_type, 16#0C#),
      997 => to_slv(opcode_type, 16#0A#),
      998 => to_slv(opcode_type, 16#06#),
      999 => to_slv(opcode_type, 16#0D#),
      1000 => to_slv(opcode_type, 16#11#),
      1001 => to_slv(opcode_type, 16#07#),
      1002 => to_slv(opcode_type, 16#04#),
      1003 => to_slv(opcode_type, 16#0F#),
      1004 => to_slv(opcode_type, 16#01#),
      1005 => to_slv(opcode_type, 16#10#),
      1006 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#05#),
      1025 => to_slv(opcode_type, 16#06#),
      1026 => to_slv(opcode_type, 16#09#),
      1027 => to_slv(opcode_type, 16#09#),
      1028 => to_slv(opcode_type, 16#0E#),
      1029 => to_slv(opcode_type, 16#0B#),
      1030 => to_slv(opcode_type, 16#06#),
      1031 => to_slv(opcode_type, 16#0E#),
      1032 => to_slv(opcode_type, 16#0D#),
      1033 => to_slv(opcode_type, 16#09#),
      1034 => to_slv(opcode_type, 16#07#),
      1035 => to_slv(opcode_type, 16#0B#),
      1036 => to_slv(opcode_type, 16#0D#),
      1037 => to_slv(opcode_type, 16#0C#),
      1038 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#09#),
      1057 => to_slv(opcode_type, 16#04#),
      1058 => to_slv(opcode_type, 16#04#),
      1059 => to_slv(opcode_type, 16#07#),
      1060 => to_slv(opcode_type, 16#0F#),
      1061 => to_slv(opcode_type, 16#0D#),
      1062 => to_slv(opcode_type, 16#01#),
      1063 => to_slv(opcode_type, 16#07#),
      1064 => to_slv(opcode_type, 16#09#),
      1065 => to_slv(opcode_type, 16#0A#),
      1066 => to_slv(opcode_type, 16#0C#),
      1067 => to_slv(opcode_type, 16#08#),
      1068 => to_slv(opcode_type, 16#0A#),
      1069 => to_slv(opcode_type, 16#0B#),
      1070 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#07#),
      1089 => to_slv(opcode_type, 16#04#),
      1090 => to_slv(opcode_type, 16#05#),
      1091 => to_slv(opcode_type, 16#06#),
      1092 => to_slv(opcode_type, 16#A0#),
      1093 => to_slv(opcode_type, 16#0B#),
      1094 => to_slv(opcode_type, 16#01#),
      1095 => to_slv(opcode_type, 16#09#),
      1096 => to_slv(opcode_type, 16#07#),
      1097 => to_slv(opcode_type, 16#0B#),
      1098 => to_slv(opcode_type, 16#0C#),
      1099 => to_slv(opcode_type, 16#09#),
      1100 => to_slv(opcode_type, 16#10#),
      1101 => to_slv(opcode_type, 16#0D#),
      1102 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#03#),
      1121 => to_slv(opcode_type, 16#07#),
      1122 => to_slv(opcode_type, 16#06#),
      1123 => to_slv(opcode_type, 16#09#),
      1124 => to_slv(opcode_type, 16#B8#),
      1125 => to_slv(opcode_type, 16#0E#),
      1126 => to_slv(opcode_type, 16#07#),
      1127 => to_slv(opcode_type, 16#0D#),
      1128 => to_slv(opcode_type, 16#0B#),
      1129 => to_slv(opcode_type, 16#07#),
      1130 => to_slv(opcode_type, 16#03#),
      1131 => to_slv(opcode_type, 16#0F#),
      1132 => to_slv(opcode_type, 16#02#),
      1133 => to_slv(opcode_type, 16#0E#),
      1134 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#02#),
      1153 => to_slv(opcode_type, 16#09#),
      1154 => to_slv(opcode_type, 16#06#),
      1155 => to_slv(opcode_type, 16#05#),
      1156 => to_slv(opcode_type, 16#0F#),
      1157 => to_slv(opcode_type, 16#02#),
      1158 => to_slv(opcode_type, 16#0C#),
      1159 => to_slv(opcode_type, 16#09#),
      1160 => to_slv(opcode_type, 16#08#),
      1161 => to_slv(opcode_type, 16#0A#),
      1162 => to_slv(opcode_type, 16#0A#),
      1163 => to_slv(opcode_type, 16#09#),
      1164 => to_slv(opcode_type, 16#0B#),
      1165 => to_slv(opcode_type, 16#10#),
      1166 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#06#),
      1185 => to_slv(opcode_type, 16#08#),
      1186 => to_slv(opcode_type, 16#05#),
      1187 => to_slv(opcode_type, 16#02#),
      1188 => to_slv(opcode_type, 16#0C#),
      1189 => to_slv(opcode_type, 16#02#),
      1190 => to_slv(opcode_type, 16#07#),
      1191 => to_slv(opcode_type, 16#10#),
      1192 => to_slv(opcode_type, 16#E1#),
      1193 => to_slv(opcode_type, 16#05#),
      1194 => to_slv(opcode_type, 16#02#),
      1195 => to_slv(opcode_type, 16#08#),
      1196 => to_slv(opcode_type, 16#0B#),
      1197 => to_slv(opcode_type, 16#0E#),
      1198 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#08#),
      1217 => to_slv(opcode_type, 16#02#),
      1218 => to_slv(opcode_type, 16#09#),
      1219 => to_slv(opcode_type, 16#09#),
      1220 => to_slv(opcode_type, 16#0B#),
      1221 => to_slv(opcode_type, 16#0D#),
      1222 => to_slv(opcode_type, 16#07#),
      1223 => to_slv(opcode_type, 16#11#),
      1224 => to_slv(opcode_type, 16#0E#),
      1225 => to_slv(opcode_type, 16#02#),
      1226 => to_slv(opcode_type, 16#02#),
      1227 => to_slv(opcode_type, 16#06#),
      1228 => to_slv(opcode_type, 16#0E#),
      1229 => to_slv(opcode_type, 16#0A#),
      1230 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#02#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#06#),
      1251 => to_slv(opcode_type, 16#04#),
      1252 => to_slv(opcode_type, 16#0B#),
      1253 => to_slv(opcode_type, 16#01#),
      1254 => to_slv(opcode_type, 16#0F#),
      1255 => to_slv(opcode_type, 16#08#),
      1256 => to_slv(opcode_type, 16#06#),
      1257 => to_slv(opcode_type, 16#0F#),
      1258 => to_slv(opcode_type, 16#11#),
      1259 => to_slv(opcode_type, 16#07#),
      1260 => to_slv(opcode_type, 16#0E#),
      1261 => to_slv(opcode_type, 16#0D#),
      1262 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#04#),
      1281 => to_slv(opcode_type, 16#07#),
      1282 => to_slv(opcode_type, 16#06#),
      1283 => to_slv(opcode_type, 16#09#),
      1284 => to_slv(opcode_type, 16#10#),
      1285 => to_slv(opcode_type, 16#10#),
      1286 => to_slv(opcode_type, 16#03#),
      1287 => to_slv(opcode_type, 16#0A#),
      1288 => to_slv(opcode_type, 16#08#),
      1289 => to_slv(opcode_type, 16#02#),
      1290 => to_slv(opcode_type, 16#11#),
      1291 => to_slv(opcode_type, 16#07#),
      1292 => to_slv(opcode_type, 16#0A#),
      1293 => to_slv(opcode_type, 16#0D#),
      1294 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#06#),
      1313 => to_slv(opcode_type, 16#07#),
      1314 => to_slv(opcode_type, 16#04#),
      1315 => to_slv(opcode_type, 16#04#),
      1316 => to_slv(opcode_type, 16#11#),
      1317 => to_slv(opcode_type, 16#08#),
      1318 => to_slv(opcode_type, 16#09#),
      1319 => to_slv(opcode_type, 16#0B#),
      1320 => to_slv(opcode_type, 16#0B#),
      1321 => to_slv(opcode_type, 16#03#),
      1322 => to_slv(opcode_type, 16#0D#),
      1323 => to_slv(opcode_type, 16#03#),
      1324 => to_slv(opcode_type, 16#05#),
      1325 => to_slv(opcode_type, 16#11#),
      1326 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#05#),
      1345 => to_slv(opcode_type, 16#06#),
      1346 => to_slv(opcode_type, 16#08#),
      1347 => to_slv(opcode_type, 16#09#),
      1348 => to_slv(opcode_type, 16#10#),
      1349 => to_slv(opcode_type, 16#D8#),
      1350 => to_slv(opcode_type, 16#04#),
      1351 => to_slv(opcode_type, 16#10#),
      1352 => to_slv(opcode_type, 16#06#),
      1353 => to_slv(opcode_type, 16#04#),
      1354 => to_slv(opcode_type, 16#0F#),
      1355 => to_slv(opcode_type, 16#07#),
      1356 => to_slv(opcode_type, 16#0E#),
      1357 => to_slv(opcode_type, 16#0B#),
      1358 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#07#),
      1377 => to_slv(opcode_type, 16#07#),
      1378 => to_slv(opcode_type, 16#01#),
      1379 => to_slv(opcode_type, 16#02#),
      1380 => to_slv(opcode_type, 16#0A#),
      1381 => to_slv(opcode_type, 16#09#),
      1382 => to_slv(opcode_type, 16#06#),
      1383 => to_slv(opcode_type, 16#0E#),
      1384 => to_slv(opcode_type, 16#0E#),
      1385 => to_slv(opcode_type, 16#06#),
      1386 => to_slv(opcode_type, 16#0D#),
      1387 => to_slv(opcode_type, 16#10#),
      1388 => to_slv(opcode_type, 16#02#),
      1389 => to_slv(opcode_type, 16#46#),
      1390 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#03#),
      1410 => to_slv(opcode_type, 16#05#),
      1411 => to_slv(opcode_type, 16#09#),
      1412 => to_slv(opcode_type, 16#83#),
      1413 => to_slv(opcode_type, 16#11#),
      1414 => to_slv(opcode_type, 16#05#),
      1415 => to_slv(opcode_type, 16#08#),
      1416 => to_slv(opcode_type, 16#06#),
      1417 => to_slv(opcode_type, 16#0E#),
      1418 => to_slv(opcode_type, 16#0D#),
      1419 => to_slv(opcode_type, 16#06#),
      1420 => to_slv(opcode_type, 16#0D#),
      1421 => to_slv(opcode_type, 16#11#),
      1422 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#08#),
      1441 => to_slv(opcode_type, 16#01#),
      1442 => to_slv(opcode_type, 16#07#),
      1443 => to_slv(opcode_type, 16#08#),
      1444 => to_slv(opcode_type, 16#0F#),
      1445 => to_slv(opcode_type, 16#0A#),
      1446 => to_slv(opcode_type, 16#04#),
      1447 => to_slv(opcode_type, 16#10#),
      1448 => to_slv(opcode_type, 16#01#),
      1449 => to_slv(opcode_type, 16#07#),
      1450 => to_slv(opcode_type, 16#08#),
      1451 => to_slv(opcode_type, 16#0E#),
      1452 => to_slv(opcode_type, 16#11#),
      1453 => to_slv(opcode_type, 16#0D#),
      1454 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#01#),
      1473 => to_slv(opcode_type, 16#06#),
      1474 => to_slv(opcode_type, 16#08#),
      1475 => to_slv(opcode_type, 16#03#),
      1476 => to_slv(opcode_type, 16#10#),
      1477 => to_slv(opcode_type, 16#03#),
      1478 => to_slv(opcode_type, 16#E9#),
      1479 => to_slv(opcode_type, 16#08#),
      1480 => to_slv(opcode_type, 16#08#),
      1481 => to_slv(opcode_type, 16#0C#),
      1482 => to_slv(opcode_type, 16#0D#),
      1483 => to_slv(opcode_type, 16#09#),
      1484 => to_slv(opcode_type, 16#0A#),
      1485 => to_slv(opcode_type, 16#0A#),
      1486 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#05#),
      1505 => to_slv(opcode_type, 16#06#),
      1506 => to_slv(opcode_type, 16#08#),
      1507 => to_slv(opcode_type, 16#07#),
      1508 => to_slv(opcode_type, 16#11#),
      1509 => to_slv(opcode_type, 16#0A#),
      1510 => to_slv(opcode_type, 16#06#),
      1511 => to_slv(opcode_type, 16#48#),
      1512 => to_slv(opcode_type, 16#11#),
      1513 => to_slv(opcode_type, 16#09#),
      1514 => to_slv(opcode_type, 16#09#),
      1515 => to_slv(opcode_type, 16#10#),
      1516 => to_slv(opcode_type, 16#0D#),
      1517 => to_slv(opcode_type, 16#0E#),
      1518 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#04#),
      1537 => to_slv(opcode_type, 16#07#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#07#),
      1540 => to_slv(opcode_type, 16#0B#),
      1541 => to_slv(opcode_type, 16#0B#),
      1542 => to_slv(opcode_type, 16#04#),
      1543 => to_slv(opcode_type, 16#0A#),
      1544 => to_slv(opcode_type, 16#07#),
      1545 => to_slv(opcode_type, 16#03#),
      1546 => to_slv(opcode_type, 16#10#),
      1547 => to_slv(opcode_type, 16#09#),
      1548 => to_slv(opcode_type, 16#10#),
      1549 => to_slv(opcode_type, 16#10#),
      1550 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#08#),
      1569 => to_slv(opcode_type, 16#05#),
      1570 => to_slv(opcode_type, 16#05#),
      1571 => to_slv(opcode_type, 16#02#),
      1572 => to_slv(opcode_type, 16#0A#),
      1573 => to_slv(opcode_type, 16#07#),
      1574 => to_slv(opcode_type, 16#01#),
      1575 => to_slv(opcode_type, 16#06#),
      1576 => to_slv(opcode_type, 16#0E#),
      1577 => to_slv(opcode_type, 16#0E#),
      1578 => to_slv(opcode_type, 16#01#),
      1579 => to_slv(opcode_type, 16#09#),
      1580 => to_slv(opcode_type, 16#0C#),
      1581 => to_slv(opcode_type, 16#11#),
      1582 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#07#),
      1601 => to_slv(opcode_type, 16#02#),
      1602 => to_slv(opcode_type, 16#02#),
      1603 => to_slv(opcode_type, 16#01#),
      1604 => to_slv(opcode_type, 16#EF#),
      1605 => to_slv(opcode_type, 16#09#),
      1606 => to_slv(opcode_type, 16#04#),
      1607 => to_slv(opcode_type, 16#08#),
      1608 => to_slv(opcode_type, 16#0D#),
      1609 => to_slv(opcode_type, 16#0A#),
      1610 => to_slv(opcode_type, 16#06#),
      1611 => to_slv(opcode_type, 16#04#),
      1612 => to_slv(opcode_type, 16#10#),
      1613 => to_slv(opcode_type, 16#11#),
      1614 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#09#),
      1633 => to_slv(opcode_type, 16#06#),
      1634 => to_slv(opcode_type, 16#04#),
      1635 => to_slv(opcode_type, 16#01#),
      1636 => to_slv(opcode_type, 16#0A#),
      1637 => to_slv(opcode_type, 16#07#),
      1638 => to_slv(opcode_type, 16#02#),
      1639 => to_slv(opcode_type, 16#0B#),
      1640 => to_slv(opcode_type, 16#04#),
      1641 => to_slv(opcode_type, 16#C8#),
      1642 => to_slv(opcode_type, 16#07#),
      1643 => to_slv(opcode_type, 16#05#),
      1644 => to_slv(opcode_type, 16#0B#),
      1645 => to_slv(opcode_type, 16#0B#),
      1646 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#07#),
      1666 => to_slv(opcode_type, 16#07#),
      1667 => to_slv(opcode_type, 16#06#),
      1668 => to_slv(opcode_type, 16#34#),
      1669 => to_slv(opcode_type, 16#0C#),
      1670 => to_slv(opcode_type, 16#03#),
      1671 => to_slv(opcode_type, 16#0E#),
      1672 => to_slv(opcode_type, 16#04#),
      1673 => to_slv(opcode_type, 16#03#),
      1674 => to_slv(opcode_type, 16#0E#),
      1675 => to_slv(opcode_type, 16#02#),
      1676 => to_slv(opcode_type, 16#01#),
      1677 => to_slv(opcode_type, 16#0F#),
      1678 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#05#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#06#),
      1699 => to_slv(opcode_type, 16#06#),
      1700 => to_slv(opcode_type, 16#C1#),
      1701 => to_slv(opcode_type, 16#0A#),
      1702 => to_slv(opcode_type, 16#04#),
      1703 => to_slv(opcode_type, 16#D8#),
      1704 => to_slv(opcode_type, 16#06#),
      1705 => to_slv(opcode_type, 16#08#),
      1706 => to_slv(opcode_type, 16#0A#),
      1707 => to_slv(opcode_type, 16#11#),
      1708 => to_slv(opcode_type, 16#03#),
      1709 => to_slv(opcode_type, 16#0A#),
      1710 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#09#),
      1729 => to_slv(opcode_type, 16#05#),
      1730 => to_slv(opcode_type, 16#08#),
      1731 => to_slv(opcode_type, 16#03#),
      1732 => to_slv(opcode_type, 16#0B#),
      1733 => to_slv(opcode_type, 16#02#),
      1734 => to_slv(opcode_type, 16#0B#),
      1735 => to_slv(opcode_type, 16#05#),
      1736 => to_slv(opcode_type, 16#08#),
      1737 => to_slv(opcode_type, 16#08#),
      1738 => to_slv(opcode_type, 16#10#),
      1739 => to_slv(opcode_type, 16#0C#),
      1740 => to_slv(opcode_type, 16#03#),
      1741 => to_slv(opcode_type, 16#0D#),
      1742 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#01#),
      1761 => to_slv(opcode_type, 16#07#),
      1762 => to_slv(opcode_type, 16#07#),
      1763 => to_slv(opcode_type, 16#09#),
      1764 => to_slv(opcode_type, 16#10#),
      1765 => to_slv(opcode_type, 16#0C#),
      1766 => to_slv(opcode_type, 16#09#),
      1767 => to_slv(opcode_type, 16#11#),
      1768 => to_slv(opcode_type, 16#10#),
      1769 => to_slv(opcode_type, 16#08#),
      1770 => to_slv(opcode_type, 16#01#),
      1771 => to_slv(opcode_type, 16#11#),
      1772 => to_slv(opcode_type, 16#03#),
      1773 => to_slv(opcode_type, 16#0D#),
      1774 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#09#),
      1793 => to_slv(opcode_type, 16#06#),
      1794 => to_slv(opcode_type, 16#09#),
      1795 => to_slv(opcode_type, 16#09#),
      1796 => to_slv(opcode_type, 16#A2#),
      1797 => to_slv(opcode_type, 16#10#),
      1798 => to_slv(opcode_type, 16#06#),
      1799 => to_slv(opcode_type, 16#0F#),
      1800 => to_slv(opcode_type, 16#0E#),
      1801 => to_slv(opcode_type, 16#04#),
      1802 => to_slv(opcode_type, 16#01#),
      1803 => to_slv(opcode_type, 16#0E#),
      1804 => to_slv(opcode_type, 16#01#),
      1805 => to_slv(opcode_type, 16#0E#),
      1806 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#06#),
      1825 => to_slv(opcode_type, 16#03#),
      1826 => to_slv(opcode_type, 16#08#),
      1827 => to_slv(opcode_type, 16#09#),
      1828 => to_slv(opcode_type, 16#0C#),
      1829 => to_slv(opcode_type, 16#2B#),
      1830 => to_slv(opcode_type, 16#05#),
      1831 => to_slv(opcode_type, 16#0C#),
      1832 => to_slv(opcode_type, 16#09#),
      1833 => to_slv(opcode_type, 16#05#),
      1834 => to_slv(opcode_type, 16#09#),
      1835 => to_slv(opcode_type, 16#0D#),
      1836 => to_slv(opcode_type, 16#0B#),
      1837 => to_slv(opcode_type, 16#5B#),
      1838 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#07#),
      1857 => to_slv(opcode_type, 16#07#),
      1858 => to_slv(opcode_type, 16#09#),
      1859 => to_slv(opcode_type, 16#04#),
      1860 => to_slv(opcode_type, 16#0D#),
      1861 => to_slv(opcode_type, 16#05#),
      1862 => to_slv(opcode_type, 16#0C#),
      1863 => to_slv(opcode_type, 16#03#),
      1864 => to_slv(opcode_type, 16#09#),
      1865 => to_slv(opcode_type, 16#0D#),
      1866 => to_slv(opcode_type, 16#0A#),
      1867 => to_slv(opcode_type, 16#06#),
      1868 => to_slv(opcode_type, 16#0E#),
      1869 => to_slv(opcode_type, 16#0E#),
      1870 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#05#),
      1889 => to_slv(opcode_type, 16#06#),
      1890 => to_slv(opcode_type, 16#09#),
      1891 => to_slv(opcode_type, 16#04#),
      1892 => to_slv(opcode_type, 16#11#),
      1893 => to_slv(opcode_type, 16#07#),
      1894 => to_slv(opcode_type, 16#0F#),
      1895 => to_slv(opcode_type, 16#0C#),
      1896 => to_slv(opcode_type, 16#06#),
      1897 => to_slv(opcode_type, 16#03#),
      1898 => to_slv(opcode_type, 16#10#),
      1899 => to_slv(opcode_type, 16#07#),
      1900 => to_slv(opcode_type, 16#11#),
      1901 => to_slv(opcode_type, 16#11#),
      1902 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#05#),
      1921 => to_slv(opcode_type, 16#07#),
      1922 => to_slv(opcode_type, 16#09#),
      1923 => to_slv(opcode_type, 16#09#),
      1924 => to_slv(opcode_type, 16#0C#),
      1925 => to_slv(opcode_type, 16#0D#),
      1926 => to_slv(opcode_type, 16#01#),
      1927 => to_slv(opcode_type, 16#0D#),
      1928 => to_slv(opcode_type, 16#06#),
      1929 => to_slv(opcode_type, 16#07#),
      1930 => to_slv(opcode_type, 16#0A#),
      1931 => to_slv(opcode_type, 16#0D#),
      1932 => to_slv(opcode_type, 16#04#),
      1933 => to_slv(opcode_type, 16#0F#),
      1934 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#03#),
      1953 => to_slv(opcode_type, 16#07#),
      1954 => to_slv(opcode_type, 16#08#),
      1955 => to_slv(opcode_type, 16#09#),
      1956 => to_slv(opcode_type, 16#11#),
      1957 => to_slv(opcode_type, 16#11#),
      1958 => to_slv(opcode_type, 16#07#),
      1959 => to_slv(opcode_type, 16#0B#),
      1960 => to_slv(opcode_type, 16#E4#),
      1961 => to_slv(opcode_type, 16#07#),
      1962 => to_slv(opcode_type, 16#06#),
      1963 => to_slv(opcode_type, 16#8E#),
      1964 => to_slv(opcode_type, 16#10#),
      1965 => to_slv(opcode_type, 16#0E#),
      1966 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#03#),
      1985 => to_slv(opcode_type, 16#07#),
      1986 => to_slv(opcode_type, 16#08#),
      1987 => to_slv(opcode_type, 16#04#),
      1988 => to_slv(opcode_type, 16#10#),
      1989 => to_slv(opcode_type, 16#08#),
      1990 => to_slv(opcode_type, 16#0F#),
      1991 => to_slv(opcode_type, 16#0A#),
      1992 => to_slv(opcode_type, 16#07#),
      1993 => to_slv(opcode_type, 16#02#),
      1994 => to_slv(opcode_type, 16#0F#),
      1995 => to_slv(opcode_type, 16#09#),
      1996 => to_slv(opcode_type, 16#8D#),
      1997 => to_slv(opcode_type, 16#0A#),
      1998 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#06#),
      2017 => to_slv(opcode_type, 16#06#),
      2018 => to_slv(opcode_type, 16#01#),
      2019 => to_slv(opcode_type, 16#06#),
      2020 => to_slv(opcode_type, 16#0D#),
      2021 => to_slv(opcode_type, 16#0F#),
      2022 => to_slv(opcode_type, 16#07#),
      2023 => to_slv(opcode_type, 16#02#),
      2024 => to_slv(opcode_type, 16#0C#),
      2025 => to_slv(opcode_type, 16#04#),
      2026 => to_slv(opcode_type, 16#0E#),
      2027 => to_slv(opcode_type, 16#08#),
      2028 => to_slv(opcode_type, 16#0C#),
      2029 => to_slv(opcode_type, 16#0F#),
      2030 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#03#),
      2049 => to_slv(opcode_type, 16#08#),
      2050 => to_slv(opcode_type, 16#08#),
      2051 => to_slv(opcode_type, 16#04#),
      2052 => to_slv(opcode_type, 16#0A#),
      2053 => to_slv(opcode_type, 16#01#),
      2054 => to_slv(opcode_type, 16#10#),
      2055 => to_slv(opcode_type, 16#07#),
      2056 => to_slv(opcode_type, 16#08#),
      2057 => to_slv(opcode_type, 16#0E#),
      2058 => to_slv(opcode_type, 16#0D#),
      2059 => to_slv(opcode_type, 16#08#),
      2060 => to_slv(opcode_type, 16#11#),
      2061 => to_slv(opcode_type, 16#0E#),
      2062 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#02#),
      2081 => to_slv(opcode_type, 16#07#),
      2082 => to_slv(opcode_type, 16#06#),
      2083 => to_slv(opcode_type, 16#09#),
      2084 => to_slv(opcode_type, 16#0A#),
      2085 => to_slv(opcode_type, 16#0A#),
      2086 => to_slv(opcode_type, 16#07#),
      2087 => to_slv(opcode_type, 16#0F#),
      2088 => to_slv(opcode_type, 16#0C#),
      2089 => to_slv(opcode_type, 16#06#),
      2090 => to_slv(opcode_type, 16#07#),
      2091 => to_slv(opcode_type, 16#10#),
      2092 => to_slv(opcode_type, 16#0C#),
      2093 => to_slv(opcode_type, 16#0A#),
      2094 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#08#),
      2113 => to_slv(opcode_type, 16#03#),
      2114 => to_slv(opcode_type, 16#07#),
      2115 => to_slv(opcode_type, 16#06#),
      2116 => to_slv(opcode_type, 16#0D#),
      2117 => to_slv(opcode_type, 16#0A#),
      2118 => to_slv(opcode_type, 16#09#),
      2119 => to_slv(opcode_type, 16#11#),
      2120 => to_slv(opcode_type, 16#10#),
      2121 => to_slv(opcode_type, 16#04#),
      2122 => to_slv(opcode_type, 16#04#),
      2123 => to_slv(opcode_type, 16#09#),
      2124 => to_slv(opcode_type, 16#0B#),
      2125 => to_slv(opcode_type, 16#92#),
      2126 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#01#),
      2145 => to_slv(opcode_type, 16#07#),
      2146 => to_slv(opcode_type, 16#06#),
      2147 => to_slv(opcode_type, 16#04#),
      2148 => to_slv(opcode_type, 16#0A#),
      2149 => to_slv(opcode_type, 16#02#),
      2150 => to_slv(opcode_type, 16#0D#),
      2151 => to_slv(opcode_type, 16#09#),
      2152 => to_slv(opcode_type, 16#09#),
      2153 => to_slv(opcode_type, 16#0A#),
      2154 => to_slv(opcode_type, 16#10#),
      2155 => to_slv(opcode_type, 16#07#),
      2156 => to_slv(opcode_type, 16#10#),
      2157 => to_slv(opcode_type, 16#0C#),
      2158 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#04#),
      2177 => to_slv(opcode_type, 16#08#),
      2178 => to_slv(opcode_type, 16#07#),
      2179 => to_slv(opcode_type, 16#07#),
      2180 => to_slv(opcode_type, 16#0D#),
      2181 => to_slv(opcode_type, 16#11#),
      2182 => to_slv(opcode_type, 16#01#),
      2183 => to_slv(opcode_type, 16#0E#),
      2184 => to_slv(opcode_type, 16#08#),
      2185 => to_slv(opcode_type, 16#02#),
      2186 => to_slv(opcode_type, 16#0E#),
      2187 => to_slv(opcode_type, 16#06#),
      2188 => to_slv(opcode_type, 16#0D#),
      2189 => to_slv(opcode_type, 16#90#),
      2190 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#01#),
      2209 => to_slv(opcode_type, 16#08#),
      2210 => to_slv(opcode_type, 16#06#),
      2211 => to_slv(opcode_type, 16#09#),
      2212 => to_slv(opcode_type, 16#0A#),
      2213 => to_slv(opcode_type, 16#11#),
      2214 => to_slv(opcode_type, 16#04#),
      2215 => to_slv(opcode_type, 16#0F#),
      2216 => to_slv(opcode_type, 16#08#),
      2217 => to_slv(opcode_type, 16#02#),
      2218 => to_slv(opcode_type, 16#2A#),
      2219 => to_slv(opcode_type, 16#07#),
      2220 => to_slv(opcode_type, 16#0D#),
      2221 => to_slv(opcode_type, 16#0B#),
      2222 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#09#),
      2241 => to_slv(opcode_type, 16#01#),
      2242 => to_slv(opcode_type, 16#02#),
      2243 => to_slv(opcode_type, 16#08#),
      2244 => to_slv(opcode_type, 16#0F#),
      2245 => to_slv(opcode_type, 16#0F#),
      2246 => to_slv(opcode_type, 16#07#),
      2247 => to_slv(opcode_type, 16#03#),
      2248 => to_slv(opcode_type, 16#05#),
      2249 => to_slv(opcode_type, 16#0D#),
      2250 => to_slv(opcode_type, 16#09#),
      2251 => to_slv(opcode_type, 16#01#),
      2252 => to_slv(opcode_type, 16#10#),
      2253 => to_slv(opcode_type, 16#11#),
      2254 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#05#),
      2273 => to_slv(opcode_type, 16#06#),
      2274 => to_slv(opcode_type, 16#06#),
      2275 => to_slv(opcode_type, 16#08#),
      2276 => to_slv(opcode_type, 16#0A#),
      2277 => to_slv(opcode_type, 16#0C#),
      2278 => to_slv(opcode_type, 16#09#),
      2279 => to_slv(opcode_type, 16#0D#),
      2280 => to_slv(opcode_type, 16#10#),
      2281 => to_slv(opcode_type, 16#06#),
      2282 => to_slv(opcode_type, 16#06#),
      2283 => to_slv(opcode_type, 16#10#),
      2284 => to_slv(opcode_type, 16#0B#),
      2285 => to_slv(opcode_type, 16#0A#),
      2286 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#01#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#06#),
      2307 => to_slv(opcode_type, 16#07#),
      2308 => to_slv(opcode_type, 16#0B#),
      2309 => to_slv(opcode_type, 16#0E#),
      2310 => to_slv(opcode_type, 16#01#),
      2311 => to_slv(opcode_type, 16#0D#),
      2312 => to_slv(opcode_type, 16#07#),
      2313 => to_slv(opcode_type, 16#03#),
      2314 => to_slv(opcode_type, 16#10#),
      2315 => to_slv(opcode_type, 16#07#),
      2316 => to_slv(opcode_type, 16#0A#),
      2317 => to_slv(opcode_type, 16#E1#),
      2318 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#01#),
      2337 => to_slv(opcode_type, 16#06#),
      2338 => to_slv(opcode_type, 16#07#),
      2339 => to_slv(opcode_type, 16#03#),
      2340 => to_slv(opcode_type, 16#0E#),
      2341 => to_slv(opcode_type, 16#01#),
      2342 => to_slv(opcode_type, 16#EA#),
      2343 => to_slv(opcode_type, 16#07#),
      2344 => to_slv(opcode_type, 16#09#),
      2345 => to_slv(opcode_type, 16#11#),
      2346 => to_slv(opcode_type, 16#0C#),
      2347 => to_slv(opcode_type, 16#07#),
      2348 => to_slv(opcode_type, 16#0F#),
      2349 => to_slv(opcode_type, 16#0F#),
      2350 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#01#),
      2369 => to_slv(opcode_type, 16#09#),
      2370 => to_slv(opcode_type, 16#09#),
      2371 => to_slv(opcode_type, 16#09#),
      2372 => to_slv(opcode_type, 16#11#),
      2373 => to_slv(opcode_type, 16#0A#),
      2374 => to_slv(opcode_type, 16#01#),
      2375 => to_slv(opcode_type, 16#0B#),
      2376 => to_slv(opcode_type, 16#08#),
      2377 => to_slv(opcode_type, 16#08#),
      2378 => to_slv(opcode_type, 16#0D#),
      2379 => to_slv(opcode_type, 16#0A#),
      2380 => to_slv(opcode_type, 16#03#),
      2381 => to_slv(opcode_type, 16#11#),
      2382 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#05#),
      2401 => to_slv(opcode_type, 16#09#),
      2402 => to_slv(opcode_type, 16#09#),
      2403 => to_slv(opcode_type, 16#05#),
      2404 => to_slv(opcode_type, 16#10#),
      2405 => to_slv(opcode_type, 16#05#),
      2406 => to_slv(opcode_type, 16#10#),
      2407 => to_slv(opcode_type, 16#09#),
      2408 => to_slv(opcode_type, 16#09#),
      2409 => to_slv(opcode_type, 16#0D#),
      2410 => to_slv(opcode_type, 16#0D#),
      2411 => to_slv(opcode_type, 16#09#),
      2412 => to_slv(opcode_type, 16#0D#),
      2413 => to_slv(opcode_type, 16#0F#),
      2414 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#02#),
      2433 => to_slv(opcode_type, 16#09#),
      2434 => to_slv(opcode_type, 16#07#),
      2435 => to_slv(opcode_type, 16#07#),
      2436 => to_slv(opcode_type, 16#0A#),
      2437 => to_slv(opcode_type, 16#0D#),
      2438 => to_slv(opcode_type, 16#04#),
      2439 => to_slv(opcode_type, 16#0E#),
      2440 => to_slv(opcode_type, 16#07#),
      2441 => to_slv(opcode_type, 16#04#),
      2442 => to_slv(opcode_type, 16#0A#),
      2443 => to_slv(opcode_type, 16#09#),
      2444 => to_slv(opcode_type, 16#0C#),
      2445 => to_slv(opcode_type, 16#0E#),
      2446 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#02#),
      2465 => to_slv(opcode_type, 16#06#),
      2466 => to_slv(opcode_type, 16#08#),
      2467 => to_slv(opcode_type, 16#08#),
      2468 => to_slv(opcode_type, 16#A6#),
      2469 => to_slv(opcode_type, 16#10#),
      2470 => to_slv(opcode_type, 16#07#),
      2471 => to_slv(opcode_type, 16#0D#),
      2472 => to_slv(opcode_type, 16#0F#),
      2473 => to_slv(opcode_type, 16#06#),
      2474 => to_slv(opcode_type, 16#07#),
      2475 => to_slv(opcode_type, 16#11#),
      2476 => to_slv(opcode_type, 16#0A#),
      2477 => to_slv(opcode_type, 16#D0#),
      2478 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#06#),
      2497 => to_slv(opcode_type, 16#01#),
      2498 => to_slv(opcode_type, 16#04#),
      2499 => to_slv(opcode_type, 16#06#),
      2500 => to_slv(opcode_type, 16#0D#),
      2501 => to_slv(opcode_type, 16#0D#),
      2502 => to_slv(opcode_type, 16#05#),
      2503 => to_slv(opcode_type, 16#07#),
      2504 => to_slv(opcode_type, 16#06#),
      2505 => to_slv(opcode_type, 16#0E#),
      2506 => to_slv(opcode_type, 16#0D#),
      2507 => to_slv(opcode_type, 16#08#),
      2508 => to_slv(opcode_type, 16#0A#),
      2509 => to_slv(opcode_type, 16#0E#),
      2510 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#06#),
      2529 => to_slv(opcode_type, 16#09#),
      2530 => to_slv(opcode_type, 16#06#),
      2531 => to_slv(opcode_type, 16#06#),
      2532 => to_slv(opcode_type, 16#10#),
      2533 => to_slv(opcode_type, 16#0E#),
      2534 => to_slv(opcode_type, 16#03#),
      2535 => to_slv(opcode_type, 16#0B#),
      2536 => to_slv(opcode_type, 16#06#),
      2537 => to_slv(opcode_type, 16#04#),
      2538 => to_slv(opcode_type, 16#0F#),
      2539 => to_slv(opcode_type, 16#05#),
      2540 => to_slv(opcode_type, 16#0C#),
      2541 => to_slv(opcode_type, 16#10#),
      2542 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#05#),
      2561 => to_slv(opcode_type, 16#06#),
      2562 => to_slv(opcode_type, 16#09#),
      2563 => to_slv(opcode_type, 16#07#),
      2564 => to_slv(opcode_type, 16#0F#),
      2565 => to_slv(opcode_type, 16#0F#),
      2566 => to_slv(opcode_type, 16#06#),
      2567 => to_slv(opcode_type, 16#11#),
      2568 => to_slv(opcode_type, 16#10#),
      2569 => to_slv(opcode_type, 16#09#),
      2570 => to_slv(opcode_type, 16#03#),
      2571 => to_slv(opcode_type, 16#0A#),
      2572 => to_slv(opcode_type, 16#04#),
      2573 => to_slv(opcode_type, 16#B2#),
      2574 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#03#),
      2593 => to_slv(opcode_type, 16#08#),
      2594 => to_slv(opcode_type, 16#09#),
      2595 => to_slv(opcode_type, 16#05#),
      2596 => to_slv(opcode_type, 16#0F#),
      2597 => to_slv(opcode_type, 16#08#),
      2598 => to_slv(opcode_type, 16#0E#),
      2599 => to_slv(opcode_type, 16#10#),
      2600 => to_slv(opcode_type, 16#09#),
      2601 => to_slv(opcode_type, 16#02#),
      2602 => to_slv(opcode_type, 16#0A#),
      2603 => to_slv(opcode_type, 16#08#),
      2604 => to_slv(opcode_type, 16#10#),
      2605 => to_slv(opcode_type, 16#0B#),
      2606 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#04#),
      2625 => to_slv(opcode_type, 16#09#),
      2626 => to_slv(opcode_type, 16#06#),
      2627 => to_slv(opcode_type, 16#05#),
      2628 => to_slv(opcode_type, 16#0A#),
      2629 => to_slv(opcode_type, 16#07#),
      2630 => to_slv(opcode_type, 16#10#),
      2631 => to_slv(opcode_type, 16#0E#),
      2632 => to_slv(opcode_type, 16#07#),
      2633 => to_slv(opcode_type, 16#09#),
      2634 => to_slv(opcode_type, 16#0C#),
      2635 => to_slv(opcode_type, 16#0F#),
      2636 => to_slv(opcode_type, 16#03#),
      2637 => to_slv(opcode_type, 16#0C#),
      2638 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#05#),
      2657 => to_slv(opcode_type, 16#07#),
      2658 => to_slv(opcode_type, 16#06#),
      2659 => to_slv(opcode_type, 16#05#),
      2660 => to_slv(opcode_type, 16#0B#),
      2661 => to_slv(opcode_type, 16#09#),
      2662 => to_slv(opcode_type, 16#0A#),
      2663 => to_slv(opcode_type, 16#0F#),
      2664 => to_slv(opcode_type, 16#07#),
      2665 => to_slv(opcode_type, 16#06#),
      2666 => to_slv(opcode_type, 16#0F#),
      2667 => to_slv(opcode_type, 16#0C#),
      2668 => to_slv(opcode_type, 16#02#),
      2669 => to_slv(opcode_type, 16#0C#),
      2670 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#02#),
      2689 => to_slv(opcode_type, 16#08#),
      2690 => to_slv(opcode_type, 16#07#),
      2691 => to_slv(opcode_type, 16#03#),
      2692 => to_slv(opcode_type, 16#0E#),
      2693 => to_slv(opcode_type, 16#04#),
      2694 => to_slv(opcode_type, 16#0C#),
      2695 => to_slv(opcode_type, 16#06#),
      2696 => to_slv(opcode_type, 16#07#),
      2697 => to_slv(opcode_type, 16#0D#),
      2698 => to_slv(opcode_type, 16#10#),
      2699 => to_slv(opcode_type, 16#09#),
      2700 => to_slv(opcode_type, 16#0E#),
      2701 => to_slv(opcode_type, 16#0F#),
      2702 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#01#),
      2721 => to_slv(opcode_type, 16#08#),
      2722 => to_slv(opcode_type, 16#06#),
      2723 => to_slv(opcode_type, 16#06#),
      2724 => to_slv(opcode_type, 16#0E#),
      2725 => to_slv(opcode_type, 16#0C#),
      2726 => to_slv(opcode_type, 16#09#),
      2727 => to_slv(opcode_type, 16#0E#),
      2728 => to_slv(opcode_type, 16#10#),
      2729 => to_slv(opcode_type, 16#06#),
      2730 => to_slv(opcode_type, 16#09#),
      2731 => to_slv(opcode_type, 16#CF#),
      2732 => to_slv(opcode_type, 16#10#),
      2733 => to_slv(opcode_type, 16#11#),
      2734 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#08#),
      2753 => to_slv(opcode_type, 16#08#),
      2754 => to_slv(opcode_type, 16#03#),
      2755 => to_slv(opcode_type, 16#08#),
      2756 => to_slv(opcode_type, 16#4B#),
      2757 => to_slv(opcode_type, 16#64#),
      2758 => to_slv(opcode_type, 16#08#),
      2759 => to_slv(opcode_type, 16#07#),
      2760 => to_slv(opcode_type, 16#0C#),
      2761 => to_slv(opcode_type, 16#0B#),
      2762 => to_slv(opcode_type, 16#03#),
      2763 => to_slv(opcode_type, 16#11#),
      2764 => to_slv(opcode_type, 16#02#),
      2765 => to_slv(opcode_type, 16#0E#),
      2766 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#02#),
      2785 => to_slv(opcode_type, 16#08#),
      2786 => to_slv(opcode_type, 16#09#),
      2787 => to_slv(opcode_type, 16#07#),
      2788 => to_slv(opcode_type, 16#0D#),
      2789 => to_slv(opcode_type, 16#0E#),
      2790 => to_slv(opcode_type, 16#01#),
      2791 => to_slv(opcode_type, 16#10#),
      2792 => to_slv(opcode_type, 16#08#),
      2793 => to_slv(opcode_type, 16#02#),
      2794 => to_slv(opcode_type, 16#0D#),
      2795 => to_slv(opcode_type, 16#08#),
      2796 => to_slv(opcode_type, 16#0B#),
      2797 => to_slv(opcode_type, 16#11#),
      2798 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#07#),
      2817 => to_slv(opcode_type, 16#07#),
      2818 => to_slv(opcode_type, 16#09#),
      2819 => to_slv(opcode_type, 16#07#),
      2820 => to_slv(opcode_type, 16#0C#),
      2821 => to_slv(opcode_type, 16#0D#),
      2822 => to_slv(opcode_type, 16#03#),
      2823 => to_slv(opcode_type, 16#10#),
      2824 => to_slv(opcode_type, 16#02#),
      2825 => to_slv(opcode_type, 16#01#),
      2826 => to_slv(opcode_type, 16#10#),
      2827 => to_slv(opcode_type, 16#02#),
      2828 => to_slv(opcode_type, 16#01#),
      2829 => to_slv(opcode_type, 16#0A#),
      2830 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#04#),
      2849 => to_slv(opcode_type, 16#09#),
      2850 => to_slv(opcode_type, 16#08#),
      2851 => to_slv(opcode_type, 16#09#),
      2852 => to_slv(opcode_type, 16#0D#),
      2853 => to_slv(opcode_type, 16#ED#),
      2854 => to_slv(opcode_type, 16#08#),
      2855 => to_slv(opcode_type, 16#0B#),
      2856 => to_slv(opcode_type, 16#5D#),
      2857 => to_slv(opcode_type, 16#07#),
      2858 => to_slv(opcode_type, 16#07#),
      2859 => to_slv(opcode_type, 16#0C#),
      2860 => to_slv(opcode_type, 16#10#),
      2861 => to_slv(opcode_type, 16#0F#),
      2862 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#05#),
      2881 => to_slv(opcode_type, 16#06#),
      2882 => to_slv(opcode_type, 16#06#),
      2883 => to_slv(opcode_type, 16#07#),
      2884 => to_slv(opcode_type, 16#0A#),
      2885 => to_slv(opcode_type, 16#11#),
      2886 => to_slv(opcode_type, 16#02#),
      2887 => to_slv(opcode_type, 16#0A#),
      2888 => to_slv(opcode_type, 16#08#),
      2889 => to_slv(opcode_type, 16#07#),
      2890 => to_slv(opcode_type, 16#0B#),
      2891 => to_slv(opcode_type, 16#11#),
      2892 => to_slv(opcode_type, 16#05#),
      2893 => to_slv(opcode_type, 16#0E#),
      2894 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#07#),
      2913 => to_slv(opcode_type, 16#06#),
      2914 => to_slv(opcode_type, 16#08#),
      2915 => to_slv(opcode_type, 16#06#),
      2916 => to_slv(opcode_type, 16#0F#),
      2917 => to_slv(opcode_type, 16#0F#),
      2918 => to_slv(opcode_type, 16#08#),
      2919 => to_slv(opcode_type, 16#0F#),
      2920 => to_slv(opcode_type, 16#0F#),
      2921 => to_slv(opcode_type, 16#08#),
      2922 => to_slv(opcode_type, 16#04#),
      2923 => to_slv(opcode_type, 16#0A#),
      2924 => to_slv(opcode_type, 16#11#),
      2925 => to_slv(opcode_type, 16#0D#),
      2926 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#06#),
      2945 => to_slv(opcode_type, 16#03#),
      2946 => to_slv(opcode_type, 16#08#),
      2947 => to_slv(opcode_type, 16#08#),
      2948 => to_slv(opcode_type, 16#0C#),
      2949 => to_slv(opcode_type, 16#10#),
      2950 => to_slv(opcode_type, 16#09#),
      2951 => to_slv(opcode_type, 16#0E#),
      2952 => to_slv(opcode_type, 16#10#),
      2953 => to_slv(opcode_type, 16#04#),
      2954 => to_slv(opcode_type, 16#03#),
      2955 => to_slv(opcode_type, 16#06#),
      2956 => to_slv(opcode_type, 16#0B#),
      2957 => to_slv(opcode_type, 16#10#),
      2958 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#02#),
      2977 => to_slv(opcode_type, 16#07#),
      2978 => to_slv(opcode_type, 16#06#),
      2979 => to_slv(opcode_type, 16#01#),
      2980 => to_slv(opcode_type, 16#0F#),
      2981 => to_slv(opcode_type, 16#06#),
      2982 => to_slv(opcode_type, 16#0B#),
      2983 => to_slv(opcode_type, 16#0F#),
      2984 => to_slv(opcode_type, 16#08#),
      2985 => to_slv(opcode_type, 16#01#),
      2986 => to_slv(opcode_type, 16#B9#),
      2987 => to_slv(opcode_type, 16#08#),
      2988 => to_slv(opcode_type, 16#0C#),
      2989 => to_slv(opcode_type, 16#7A#),
      2990 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#05#),
      3009 => to_slv(opcode_type, 16#06#),
      3010 => to_slv(opcode_type, 16#09#),
      3011 => to_slv(opcode_type, 16#09#),
      3012 => to_slv(opcode_type, 16#11#),
      3013 => to_slv(opcode_type, 16#0C#),
      3014 => to_slv(opcode_type, 16#08#),
      3015 => to_slv(opcode_type, 16#0A#),
      3016 => to_slv(opcode_type, 16#10#),
      3017 => to_slv(opcode_type, 16#07#),
      3018 => to_slv(opcode_type, 16#09#),
      3019 => to_slv(opcode_type, 16#63#),
      3020 => to_slv(opcode_type, 16#0D#),
      3021 => to_slv(opcode_type, 16#10#),
      3022 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#06#),
      3041 => to_slv(opcode_type, 16#04#),
      3042 => to_slv(opcode_type, 16#02#),
      3043 => to_slv(opcode_type, 16#09#),
      3044 => to_slv(opcode_type, 16#0B#),
      3045 => to_slv(opcode_type, 16#0A#),
      3046 => to_slv(opcode_type, 16#06#),
      3047 => to_slv(opcode_type, 16#04#),
      3048 => to_slv(opcode_type, 16#08#),
      3049 => to_slv(opcode_type, 16#0E#),
      3050 => to_slv(opcode_type, 16#10#),
      3051 => to_slv(opcode_type, 16#09#),
      3052 => to_slv(opcode_type, 16#11#),
      3053 => to_slv(opcode_type, 16#0D#),
      3054 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#07#),
      3073 => to_slv(opcode_type, 16#07#),
      3074 => to_slv(opcode_type, 16#02#),
      3075 => to_slv(opcode_type, 16#03#),
      3076 => to_slv(opcode_type, 16#0F#),
      3077 => to_slv(opcode_type, 16#03#),
      3078 => to_slv(opcode_type, 16#07#),
      3079 => to_slv(opcode_type, 16#0E#),
      3080 => to_slv(opcode_type, 16#11#),
      3081 => to_slv(opcode_type, 16#06#),
      3082 => to_slv(opcode_type, 16#04#),
      3083 => to_slv(opcode_type, 16#04#),
      3084 => to_slv(opcode_type, 16#96#),
      3085 => to_slv(opcode_type, 16#0C#),
      3086 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#09#),
      3105 => to_slv(opcode_type, 16#09#),
      3106 => to_slv(opcode_type, 16#04#),
      3107 => to_slv(opcode_type, 16#04#),
      3108 => to_slv(opcode_type, 16#0F#),
      3109 => to_slv(opcode_type, 16#03#),
      3110 => to_slv(opcode_type, 16#06#),
      3111 => to_slv(opcode_type, 16#0D#),
      3112 => to_slv(opcode_type, 16#3E#),
      3113 => to_slv(opcode_type, 16#02#),
      3114 => to_slv(opcode_type, 16#05#),
      3115 => to_slv(opcode_type, 16#09#),
      3116 => to_slv(opcode_type, 16#10#),
      3117 => to_slv(opcode_type, 16#0D#),
      3118 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#08#),
      3137 => to_slv(opcode_type, 16#04#),
      3138 => to_slv(opcode_type, 16#01#),
      3139 => to_slv(opcode_type, 16#07#),
      3140 => to_slv(opcode_type, 16#0A#),
      3141 => to_slv(opcode_type, 16#0B#),
      3142 => to_slv(opcode_type, 16#01#),
      3143 => to_slv(opcode_type, 16#08#),
      3144 => to_slv(opcode_type, 16#06#),
      3145 => to_slv(opcode_type, 16#0C#),
      3146 => to_slv(opcode_type, 16#10#),
      3147 => to_slv(opcode_type, 16#06#),
      3148 => to_slv(opcode_type, 16#0C#),
      3149 => to_slv(opcode_type, 16#0E#),
      3150 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#05#),
      3169 => to_slv(opcode_type, 16#07#),
      3170 => to_slv(opcode_type, 16#08#),
      3171 => to_slv(opcode_type, 16#01#),
      3172 => to_slv(opcode_type, 16#0A#),
      3173 => to_slv(opcode_type, 16#08#),
      3174 => to_slv(opcode_type, 16#0C#),
      3175 => to_slv(opcode_type, 16#0C#),
      3176 => to_slv(opcode_type, 16#06#),
      3177 => to_slv(opcode_type, 16#06#),
      3178 => to_slv(opcode_type, 16#0B#),
      3179 => to_slv(opcode_type, 16#0D#),
      3180 => to_slv(opcode_type, 16#05#),
      3181 => to_slv(opcode_type, 16#0E#),
      3182 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#01#),
      3201 => to_slv(opcode_type, 16#09#),
      3202 => to_slv(opcode_type, 16#06#),
      3203 => to_slv(opcode_type, 16#09#),
      3204 => to_slv(opcode_type, 16#11#),
      3205 => to_slv(opcode_type, 16#0D#),
      3206 => to_slv(opcode_type, 16#09#),
      3207 => to_slv(opcode_type, 16#0C#),
      3208 => to_slv(opcode_type, 16#0E#),
      3209 => to_slv(opcode_type, 16#07#),
      3210 => to_slv(opcode_type, 16#01#),
      3211 => to_slv(opcode_type, 16#0F#),
      3212 => to_slv(opcode_type, 16#03#),
      3213 => to_slv(opcode_type, 16#79#),
      3214 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#09#),
      3233 => to_slv(opcode_type, 16#02#),
      3234 => to_slv(opcode_type, 16#05#),
      3235 => to_slv(opcode_type, 16#03#),
      3236 => to_slv(opcode_type, 16#0C#),
      3237 => to_slv(opcode_type, 16#06#),
      3238 => to_slv(opcode_type, 16#03#),
      3239 => to_slv(opcode_type, 16#04#),
      3240 => to_slv(opcode_type, 16#0F#),
      3241 => to_slv(opcode_type, 16#07#),
      3242 => to_slv(opcode_type, 16#04#),
      3243 => to_slv(opcode_type, 16#10#),
      3244 => to_slv(opcode_type, 16#03#),
      3245 => to_slv(opcode_type, 16#0A#),
      3246 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#09#),
      3265 => to_slv(opcode_type, 16#04#),
      3266 => to_slv(opcode_type, 16#09#),
      3267 => to_slv(opcode_type, 16#06#),
      3268 => to_slv(opcode_type, 16#0C#),
      3269 => to_slv(opcode_type, 16#0B#),
      3270 => to_slv(opcode_type, 16#09#),
      3271 => to_slv(opcode_type, 16#10#),
      3272 => to_slv(opcode_type, 16#B1#),
      3273 => to_slv(opcode_type, 16#03#),
      3274 => to_slv(opcode_type, 16#02#),
      3275 => to_slv(opcode_type, 16#09#),
      3276 => to_slv(opcode_type, 16#0A#),
      3277 => to_slv(opcode_type, 16#0D#),
      3278 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#02#),
      3297 => to_slv(opcode_type, 16#09#),
      3298 => to_slv(opcode_type, 16#06#),
      3299 => to_slv(opcode_type, 16#04#),
      3300 => to_slv(opcode_type, 16#0A#),
      3301 => to_slv(opcode_type, 16#03#),
      3302 => to_slv(opcode_type, 16#C9#),
      3303 => to_slv(opcode_type, 16#09#),
      3304 => to_slv(opcode_type, 16#09#),
      3305 => to_slv(opcode_type, 16#0E#),
      3306 => to_slv(opcode_type, 16#0B#),
      3307 => to_slv(opcode_type, 16#06#),
      3308 => to_slv(opcode_type, 16#0E#),
      3309 => to_slv(opcode_type, 16#10#),
      3310 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#02#),
      3329 => to_slv(opcode_type, 16#09#),
      3330 => to_slv(opcode_type, 16#07#),
      3331 => to_slv(opcode_type, 16#04#),
      3332 => to_slv(opcode_type, 16#0B#),
      3333 => to_slv(opcode_type, 16#03#),
      3334 => to_slv(opcode_type, 16#3A#),
      3335 => to_slv(opcode_type, 16#09#),
      3336 => to_slv(opcode_type, 16#07#),
      3337 => to_slv(opcode_type, 16#0E#),
      3338 => to_slv(opcode_type, 16#0F#),
      3339 => to_slv(opcode_type, 16#07#),
      3340 => to_slv(opcode_type, 16#0F#),
      3341 => to_slv(opcode_type, 16#0A#),
      3342 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#09#),
      3361 => to_slv(opcode_type, 16#03#),
      3362 => to_slv(opcode_type, 16#01#),
      3363 => to_slv(opcode_type, 16#05#),
      3364 => to_slv(opcode_type, 16#0E#),
      3365 => to_slv(opcode_type, 16#06#),
      3366 => to_slv(opcode_type, 16#09#),
      3367 => to_slv(opcode_type, 16#09#),
      3368 => to_slv(opcode_type, 16#0E#),
      3369 => to_slv(opcode_type, 16#0E#),
      3370 => to_slv(opcode_type, 16#02#),
      3371 => to_slv(opcode_type, 16#0C#),
      3372 => to_slv(opcode_type, 16#03#),
      3373 => to_slv(opcode_type, 16#10#),
      3374 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#01#),
      3393 => to_slv(opcode_type, 16#07#),
      3394 => to_slv(opcode_type, 16#09#),
      3395 => to_slv(opcode_type, 16#02#),
      3396 => to_slv(opcode_type, 16#0D#),
      3397 => to_slv(opcode_type, 16#06#),
      3398 => to_slv(opcode_type, 16#11#),
      3399 => to_slv(opcode_type, 16#ED#),
      3400 => to_slv(opcode_type, 16#06#),
      3401 => to_slv(opcode_type, 16#06#),
      3402 => to_slv(opcode_type, 16#87#),
      3403 => to_slv(opcode_type, 16#0C#),
      3404 => to_slv(opcode_type, 16#01#),
      3405 => to_slv(opcode_type, 16#62#),
      3406 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#01#),
      3425 => to_slv(opcode_type, 16#06#),
      3426 => to_slv(opcode_type, 16#06#),
      3427 => to_slv(opcode_type, 16#06#),
      3428 => to_slv(opcode_type, 16#5C#),
      3429 => to_slv(opcode_type, 16#0F#),
      3430 => to_slv(opcode_type, 16#01#),
      3431 => to_slv(opcode_type, 16#0C#),
      3432 => to_slv(opcode_type, 16#06#),
      3433 => to_slv(opcode_type, 16#04#),
      3434 => to_slv(opcode_type, 16#0E#),
      3435 => to_slv(opcode_type, 16#06#),
      3436 => to_slv(opcode_type, 16#0D#),
      3437 => to_slv(opcode_type, 16#0F#),
      3438 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#03#),
      3457 => to_slv(opcode_type, 16#09#),
      3458 => to_slv(opcode_type, 16#06#),
      3459 => to_slv(opcode_type, 16#02#),
      3460 => to_slv(opcode_type, 16#0A#),
      3461 => to_slv(opcode_type, 16#09#),
      3462 => to_slv(opcode_type, 16#0A#),
      3463 => to_slv(opcode_type, 16#0A#),
      3464 => to_slv(opcode_type, 16#08#),
      3465 => to_slv(opcode_type, 16#05#),
      3466 => to_slv(opcode_type, 16#0F#),
      3467 => to_slv(opcode_type, 16#09#),
      3468 => to_slv(opcode_type, 16#10#),
      3469 => to_slv(opcode_type, 16#0F#),
      3470 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#02#),
      3489 => to_slv(opcode_type, 16#08#),
      3490 => to_slv(opcode_type, 16#09#),
      3491 => to_slv(opcode_type, 16#04#),
      3492 => to_slv(opcode_type, 16#0B#),
      3493 => to_slv(opcode_type, 16#02#),
      3494 => to_slv(opcode_type, 16#0A#),
      3495 => to_slv(opcode_type, 16#09#),
      3496 => to_slv(opcode_type, 16#07#),
      3497 => to_slv(opcode_type, 16#75#),
      3498 => to_slv(opcode_type, 16#CB#),
      3499 => to_slv(opcode_type, 16#09#),
      3500 => to_slv(opcode_type, 16#0F#),
      3501 => to_slv(opcode_type, 16#10#),
      3502 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#04#),
      3521 => to_slv(opcode_type, 16#09#),
      3522 => to_slv(opcode_type, 16#06#),
      3523 => to_slv(opcode_type, 16#09#),
      3524 => to_slv(opcode_type, 16#11#),
      3525 => to_slv(opcode_type, 16#0D#),
      3526 => to_slv(opcode_type, 16#08#),
      3527 => to_slv(opcode_type, 16#11#),
      3528 => to_slv(opcode_type, 16#0B#),
      3529 => to_slv(opcode_type, 16#07#),
      3530 => to_slv(opcode_type, 16#04#),
      3531 => to_slv(opcode_type, 16#0E#),
      3532 => to_slv(opcode_type, 16#02#),
      3533 => to_slv(opcode_type, 16#0F#),
      3534 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#02#),
      3553 => to_slv(opcode_type, 16#07#),
      3554 => to_slv(opcode_type, 16#06#),
      3555 => to_slv(opcode_type, 16#09#),
      3556 => to_slv(opcode_type, 16#0F#),
      3557 => to_slv(opcode_type, 16#C5#),
      3558 => to_slv(opcode_type, 16#08#),
      3559 => to_slv(opcode_type, 16#0E#),
      3560 => to_slv(opcode_type, 16#0B#),
      3561 => to_slv(opcode_type, 16#08#),
      3562 => to_slv(opcode_type, 16#05#),
      3563 => to_slv(opcode_type, 16#0F#),
      3564 => to_slv(opcode_type, 16#05#),
      3565 => to_slv(opcode_type, 16#0E#),
      3566 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#01#),
      3585 => to_slv(opcode_type, 16#06#),
      3586 => to_slv(opcode_type, 16#06#),
      3587 => to_slv(opcode_type, 16#06#),
      3588 => to_slv(opcode_type, 16#0F#),
      3589 => to_slv(opcode_type, 16#50#),
      3590 => to_slv(opcode_type, 16#06#),
      3591 => to_slv(opcode_type, 16#98#),
      3592 => to_slv(opcode_type, 16#10#),
      3593 => to_slv(opcode_type, 16#09#),
      3594 => to_slv(opcode_type, 16#08#),
      3595 => to_slv(opcode_type, 16#0B#),
      3596 => to_slv(opcode_type, 16#0C#),
      3597 => to_slv(opcode_type, 16#C4#),
      3598 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#04#),
      3617 => to_slv(opcode_type, 16#07#),
      3618 => to_slv(opcode_type, 16#09#),
      3619 => to_slv(opcode_type, 16#06#),
      3620 => to_slv(opcode_type, 16#A5#),
      3621 => to_slv(opcode_type, 16#10#),
      3622 => to_slv(opcode_type, 16#01#),
      3623 => to_slv(opcode_type, 16#57#),
      3624 => to_slv(opcode_type, 16#07#),
      3625 => to_slv(opcode_type, 16#01#),
      3626 => to_slv(opcode_type, 16#0A#),
      3627 => to_slv(opcode_type, 16#09#),
      3628 => to_slv(opcode_type, 16#0B#),
      3629 => to_slv(opcode_type, 16#0A#),
      3630 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#03#),
      3649 => to_slv(opcode_type, 16#06#),
      3650 => to_slv(opcode_type, 16#06#),
      3651 => to_slv(opcode_type, 16#08#),
      3652 => to_slv(opcode_type, 16#78#),
      3653 => to_slv(opcode_type, 16#11#),
      3654 => to_slv(opcode_type, 16#07#),
      3655 => to_slv(opcode_type, 16#0E#),
      3656 => to_slv(opcode_type, 16#0B#),
      3657 => to_slv(opcode_type, 16#08#),
      3658 => to_slv(opcode_type, 16#09#),
      3659 => to_slv(opcode_type, 16#0A#),
      3660 => to_slv(opcode_type, 16#0C#),
      3661 => to_slv(opcode_type, 16#0D#),
      3662 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#08#),
      3681 => to_slv(opcode_type, 16#02#),
      3682 => to_slv(opcode_type, 16#03#),
      3683 => to_slv(opcode_type, 16#09#),
      3684 => to_slv(opcode_type, 16#F2#),
      3685 => to_slv(opcode_type, 16#0C#),
      3686 => to_slv(opcode_type, 16#04#),
      3687 => to_slv(opcode_type, 16#06#),
      3688 => to_slv(opcode_type, 16#08#),
      3689 => to_slv(opcode_type, 16#0B#),
      3690 => to_slv(opcode_type, 16#11#),
      3691 => to_slv(opcode_type, 16#06#),
      3692 => to_slv(opcode_type, 16#0E#),
      3693 => to_slv(opcode_type, 16#0F#),
      3694 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#05#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#06#),
      3715 => to_slv(opcode_type, 16#02#),
      3716 => to_slv(opcode_type, 16#0A#),
      3717 => to_slv(opcode_type, 16#08#),
      3718 => to_slv(opcode_type, 16#11#),
      3719 => to_slv(opcode_type, 16#0F#),
      3720 => to_slv(opcode_type, 16#08#),
      3721 => to_slv(opcode_type, 16#08#),
      3722 => to_slv(opcode_type, 16#0E#),
      3723 => to_slv(opcode_type, 16#0B#),
      3724 => to_slv(opcode_type, 16#01#),
      3725 => to_slv(opcode_type, 16#0C#),
      3726 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#06#),
      3745 => to_slv(opcode_type, 16#07#),
      3746 => to_slv(opcode_type, 16#06#),
      3747 => to_slv(opcode_type, 16#07#),
      3748 => to_slv(opcode_type, 16#0F#),
      3749 => to_slv(opcode_type, 16#0C#),
      3750 => to_slv(opcode_type, 16#03#),
      3751 => to_slv(opcode_type, 16#F4#),
      3752 => to_slv(opcode_type, 16#03#),
      3753 => to_slv(opcode_type, 16#08#),
      3754 => to_slv(opcode_type, 16#0F#),
      3755 => to_slv(opcode_type, 16#A4#),
      3756 => to_slv(opcode_type, 16#01#),
      3757 => to_slv(opcode_type, 16#0F#),
      3758 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#09#),
      3777 => to_slv(opcode_type, 16#07#),
      3778 => to_slv(opcode_type, 16#02#),
      3779 => to_slv(opcode_type, 16#09#),
      3780 => to_slv(opcode_type, 16#0D#),
      3781 => to_slv(opcode_type, 16#0E#),
      3782 => to_slv(opcode_type, 16#02#),
      3783 => to_slv(opcode_type, 16#03#),
      3784 => to_slv(opcode_type, 16#46#),
      3785 => to_slv(opcode_type, 16#07#),
      3786 => to_slv(opcode_type, 16#04#),
      3787 => to_slv(opcode_type, 16#01#),
      3788 => to_slv(opcode_type, 16#10#),
      3789 => to_slv(opcode_type, 16#11#),
      3790 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#09#),
      3809 => to_slv(opcode_type, 16#01#),
      3810 => to_slv(opcode_type, 16#09#),
      3811 => to_slv(opcode_type, 16#04#),
      3812 => to_slv(opcode_type, 16#45#),
      3813 => to_slv(opcode_type, 16#09#),
      3814 => to_slv(opcode_type, 16#0E#),
      3815 => to_slv(opcode_type, 16#0D#),
      3816 => to_slv(opcode_type, 16#06#),
      3817 => to_slv(opcode_type, 16#01#),
      3818 => to_slv(opcode_type, 16#02#),
      3819 => to_slv(opcode_type, 16#0F#),
      3820 => to_slv(opcode_type, 16#02#),
      3821 => to_slv(opcode_type, 16#11#),
      3822 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#03#),
      3841 => to_slv(opcode_type, 16#06#),
      3842 => to_slv(opcode_type, 16#08#),
      3843 => to_slv(opcode_type, 16#03#),
      3844 => to_slv(opcode_type, 16#0F#),
      3845 => to_slv(opcode_type, 16#04#),
      3846 => to_slv(opcode_type, 16#10#),
      3847 => to_slv(opcode_type, 16#06#),
      3848 => to_slv(opcode_type, 16#08#),
      3849 => to_slv(opcode_type, 16#0B#),
      3850 => to_slv(opcode_type, 16#0B#),
      3851 => to_slv(opcode_type, 16#09#),
      3852 => to_slv(opcode_type, 16#0C#),
      3853 => to_slv(opcode_type, 16#0B#),
      3854 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#04#),
      3873 => to_slv(opcode_type, 16#08#),
      3874 => to_slv(opcode_type, 16#09#),
      3875 => to_slv(opcode_type, 16#03#),
      3876 => to_slv(opcode_type, 16#0C#),
      3877 => to_slv(opcode_type, 16#07#),
      3878 => to_slv(opcode_type, 16#0D#),
      3879 => to_slv(opcode_type, 16#0E#),
      3880 => to_slv(opcode_type, 16#06#),
      3881 => to_slv(opcode_type, 16#03#),
      3882 => to_slv(opcode_type, 16#10#),
      3883 => to_slv(opcode_type, 16#06#),
      3884 => to_slv(opcode_type, 16#0B#),
      3885 => to_slv(opcode_type, 16#0F#),
      3886 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#03#),
      3905 => to_slv(opcode_type, 16#06#),
      3906 => to_slv(opcode_type, 16#09#),
      3907 => to_slv(opcode_type, 16#07#),
      3908 => to_slv(opcode_type, 16#0B#),
      3909 => to_slv(opcode_type, 16#10#),
      3910 => to_slv(opcode_type, 16#01#),
      3911 => to_slv(opcode_type, 16#11#),
      3912 => to_slv(opcode_type, 16#06#),
      3913 => to_slv(opcode_type, 16#01#),
      3914 => to_slv(opcode_type, 16#0C#),
      3915 => to_slv(opcode_type, 16#09#),
      3916 => to_slv(opcode_type, 16#0D#),
      3917 => to_slv(opcode_type, 16#0B#),
      3918 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#01#),
      3937 => to_slv(opcode_type, 16#07#),
      3938 => to_slv(opcode_type, 16#08#),
      3939 => to_slv(opcode_type, 16#02#),
      3940 => to_slv(opcode_type, 16#0D#),
      3941 => to_slv(opcode_type, 16#03#),
      3942 => to_slv(opcode_type, 16#0F#),
      3943 => to_slv(opcode_type, 16#08#),
      3944 => to_slv(opcode_type, 16#09#),
      3945 => to_slv(opcode_type, 16#E5#),
      3946 => to_slv(opcode_type, 16#0C#),
      3947 => to_slv(opcode_type, 16#06#),
      3948 => to_slv(opcode_type, 16#11#),
      3949 => to_slv(opcode_type, 16#0B#),
      3950 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#05#),
      3969 => to_slv(opcode_type, 16#09#),
      3970 => to_slv(opcode_type, 16#09#),
      3971 => to_slv(opcode_type, 16#01#),
      3972 => to_slv(opcode_type, 16#82#),
      3973 => to_slv(opcode_type, 16#02#),
      3974 => to_slv(opcode_type, 16#0E#),
      3975 => to_slv(opcode_type, 16#07#),
      3976 => to_slv(opcode_type, 16#07#),
      3977 => to_slv(opcode_type, 16#6D#),
      3978 => to_slv(opcode_type, 16#0F#),
      3979 => to_slv(opcode_type, 16#06#),
      3980 => to_slv(opcode_type, 16#0A#),
      3981 => to_slv(opcode_type, 16#0B#),
      3982 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#06#),
      4001 => to_slv(opcode_type, 16#03#),
      4002 => to_slv(opcode_type, 16#08#),
      4003 => to_slv(opcode_type, 16#01#),
      4004 => to_slv(opcode_type, 16#11#),
      4005 => to_slv(opcode_type, 16#07#),
      4006 => to_slv(opcode_type, 16#0C#),
      4007 => to_slv(opcode_type, 16#10#),
      4008 => to_slv(opcode_type, 16#05#),
      4009 => to_slv(opcode_type, 16#08#),
      4010 => to_slv(opcode_type, 16#02#),
      4011 => to_slv(opcode_type, 16#0B#),
      4012 => to_slv(opcode_type, 16#05#),
      4013 => to_slv(opcode_type, 16#10#),
      4014 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#01#),
      4033 => to_slv(opcode_type, 16#06#),
      4034 => to_slv(opcode_type, 16#08#),
      4035 => to_slv(opcode_type, 16#06#),
      4036 => to_slv(opcode_type, 16#0B#),
      4037 => to_slv(opcode_type, 16#0E#),
      4038 => to_slv(opcode_type, 16#09#),
      4039 => to_slv(opcode_type, 16#0E#),
      4040 => to_slv(opcode_type, 16#1A#),
      4041 => to_slv(opcode_type, 16#06#),
      4042 => to_slv(opcode_type, 16#06#),
      4043 => to_slv(opcode_type, 16#0D#),
      4044 => to_slv(opcode_type, 16#0F#),
      4045 => to_slv(opcode_type, 16#8B#),
      4046 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#09#),
      4065 => to_slv(opcode_type, 16#08#),
      4066 => to_slv(opcode_type, 16#02#),
      4067 => to_slv(opcode_type, 16#06#),
      4068 => to_slv(opcode_type, 16#0D#),
      4069 => to_slv(opcode_type, 16#0C#),
      4070 => to_slv(opcode_type, 16#02#),
      4071 => to_slv(opcode_type, 16#01#),
      4072 => to_slv(opcode_type, 16#0B#),
      4073 => to_slv(opcode_type, 16#09#),
      4074 => to_slv(opcode_type, 16#03#),
      4075 => to_slv(opcode_type, 16#04#),
      4076 => to_slv(opcode_type, 16#0D#),
      4077 => to_slv(opcode_type, 16#0D#),
      4078 to 4095 => (others => '0')
  ),

    -- Bin `15`...
    14 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#04#),
      1 => to_slv(opcode_type, 16#08#),
      2 => to_slv(opcode_type, 16#06#),
      3 => to_slv(opcode_type, 16#08#),
      4 => to_slv(opcode_type, 16#0C#),
      5 => to_slv(opcode_type, 16#0A#),
      6 => to_slv(opcode_type, 16#03#),
      7 => to_slv(opcode_type, 16#0B#),
      8 => to_slv(opcode_type, 16#08#),
      9 => to_slv(opcode_type, 16#09#),
      10 => to_slv(opcode_type, 16#C1#),
      11 => to_slv(opcode_type, 16#0B#),
      12 => to_slv(opcode_type, 16#09#),
      13 => to_slv(opcode_type, 16#0C#),
      14 => to_slv(opcode_type, 16#0A#),
      15 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#01#),
      33 => to_slv(opcode_type, 16#06#),
      34 => to_slv(opcode_type, 16#08#),
      35 => to_slv(opcode_type, 16#09#),
      36 => to_slv(opcode_type, 16#0E#),
      37 => to_slv(opcode_type, 16#10#),
      38 => to_slv(opcode_type, 16#04#),
      39 => to_slv(opcode_type, 16#0E#),
      40 => to_slv(opcode_type, 16#09#),
      41 => to_slv(opcode_type, 16#08#),
      42 => to_slv(opcode_type, 16#7B#),
      43 => to_slv(opcode_type, 16#6C#),
      44 => to_slv(opcode_type, 16#07#),
      45 => to_slv(opcode_type, 16#0F#),
      46 => to_slv(opcode_type, 16#0B#),
      47 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#06#),
      65 => to_slv(opcode_type, 16#09#),
      66 => to_slv(opcode_type, 16#04#),
      67 => to_slv(opcode_type, 16#07#),
      68 => to_slv(opcode_type, 16#0F#),
      69 => to_slv(opcode_type, 16#0B#),
      70 => to_slv(opcode_type, 16#05#),
      71 => to_slv(opcode_type, 16#09#),
      72 => to_slv(opcode_type, 16#0C#),
      73 => to_slv(opcode_type, 16#11#),
      74 => to_slv(opcode_type, 16#07#),
      75 => to_slv(opcode_type, 16#09#),
      76 => to_slv(opcode_type, 16#0D#),
      77 => to_slv(opcode_type, 16#11#),
      78 => to_slv(opcode_type, 16#10#),
      79 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#01#),
      97 => to_slv(opcode_type, 16#08#),
      98 => to_slv(opcode_type, 16#09#),
      99 => to_slv(opcode_type, 16#05#),
      100 => to_slv(opcode_type, 16#0B#),
      101 => to_slv(opcode_type, 16#08#),
      102 => to_slv(opcode_type, 16#0A#),
      103 => to_slv(opcode_type, 16#0A#),
      104 => to_slv(opcode_type, 16#07#),
      105 => to_slv(opcode_type, 16#08#),
      106 => to_slv(opcode_type, 16#0C#),
      107 => to_slv(opcode_type, 16#0C#),
      108 => to_slv(opcode_type, 16#06#),
      109 => to_slv(opcode_type, 16#0B#),
      110 => to_slv(opcode_type, 16#10#),
      111 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#05#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#07#),
      131 => to_slv(opcode_type, 16#07#),
      132 => to_slv(opcode_type, 16#0F#),
      133 => to_slv(opcode_type, 16#0B#),
      134 => to_slv(opcode_type, 16#09#),
      135 => to_slv(opcode_type, 16#0C#),
      136 => to_slv(opcode_type, 16#11#),
      137 => to_slv(opcode_type, 16#07#),
      138 => to_slv(opcode_type, 16#05#),
      139 => to_slv(opcode_type, 16#10#),
      140 => to_slv(opcode_type, 16#06#),
      141 => to_slv(opcode_type, 16#0C#),
      142 => to_slv(opcode_type, 16#0F#),
      143 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#02#),
      161 => to_slv(opcode_type, 16#09#),
      162 => to_slv(opcode_type, 16#07#),
      163 => to_slv(opcode_type, 16#07#),
      164 => to_slv(opcode_type, 16#0B#),
      165 => to_slv(opcode_type, 16#0C#),
      166 => to_slv(opcode_type, 16#09#),
      167 => to_slv(opcode_type, 16#0C#),
      168 => to_slv(opcode_type, 16#0C#),
      169 => to_slv(opcode_type, 16#08#),
      170 => to_slv(opcode_type, 16#04#),
      171 => to_slv(opcode_type, 16#59#),
      172 => to_slv(opcode_type, 16#09#),
      173 => to_slv(opcode_type, 16#0E#),
      174 => to_slv(opcode_type, 16#0B#),
      175 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#01#),
      193 => to_slv(opcode_type, 16#06#),
      194 => to_slv(opcode_type, 16#09#),
      195 => to_slv(opcode_type, 16#08#),
      196 => to_slv(opcode_type, 16#0D#),
      197 => to_slv(opcode_type, 16#0B#),
      198 => to_slv(opcode_type, 16#04#),
      199 => to_slv(opcode_type, 16#11#),
      200 => to_slv(opcode_type, 16#09#),
      201 => to_slv(opcode_type, 16#09#),
      202 => to_slv(opcode_type, 16#0D#),
      203 => to_slv(opcode_type, 16#10#),
      204 => to_slv(opcode_type, 16#07#),
      205 => to_slv(opcode_type, 16#11#),
      206 => to_slv(opcode_type, 16#A7#),
      207 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#04#),
      225 => to_slv(opcode_type, 16#08#),
      226 => to_slv(opcode_type, 16#06#),
      227 => to_slv(opcode_type, 16#04#),
      228 => to_slv(opcode_type, 16#10#),
      229 => to_slv(opcode_type, 16#07#),
      230 => to_slv(opcode_type, 16#11#),
      231 => to_slv(opcode_type, 16#0B#),
      232 => to_slv(opcode_type, 16#06#),
      233 => to_slv(opcode_type, 16#09#),
      234 => to_slv(opcode_type, 16#0F#),
      235 => to_slv(opcode_type, 16#0D#),
      236 => to_slv(opcode_type, 16#06#),
      237 => to_slv(opcode_type, 16#11#),
      238 => to_slv(opcode_type, 16#11#),
      239 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#07#),
      257 => to_slv(opcode_type, 16#09#),
      258 => to_slv(opcode_type, 16#09#),
      259 => to_slv(opcode_type, 16#06#),
      260 => to_slv(opcode_type, 16#0D#),
      261 => to_slv(opcode_type, 16#0D#),
      262 => to_slv(opcode_type, 16#08#),
      263 => to_slv(opcode_type, 16#0C#),
      264 => to_slv(opcode_type, 16#0D#),
      265 => to_slv(opcode_type, 16#02#),
      266 => to_slv(opcode_type, 16#07#),
      267 => to_slv(opcode_type, 16#0B#),
      268 => to_slv(opcode_type, 16#0E#),
      269 => to_slv(opcode_type, 16#01#),
      270 => to_slv(opcode_type, 16#0C#),
      271 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#03#),
      289 => to_slv(opcode_type, 16#07#),
      290 => to_slv(opcode_type, 16#08#),
      291 => to_slv(opcode_type, 16#05#),
      292 => to_slv(opcode_type, 16#10#),
      293 => to_slv(opcode_type, 16#08#),
      294 => to_slv(opcode_type, 16#0A#),
      295 => to_slv(opcode_type, 16#0F#),
      296 => to_slv(opcode_type, 16#07#),
      297 => to_slv(opcode_type, 16#08#),
      298 => to_slv(opcode_type, 16#0B#),
      299 => to_slv(opcode_type, 16#11#),
      300 => to_slv(opcode_type, 16#07#),
      301 => to_slv(opcode_type, 16#0B#),
      302 => to_slv(opcode_type, 16#11#),
      303 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#04#),
      321 => to_slv(opcode_type, 16#08#),
      322 => to_slv(opcode_type, 16#08#),
      323 => to_slv(opcode_type, 16#01#),
      324 => to_slv(opcode_type, 16#0D#),
      325 => to_slv(opcode_type, 16#09#),
      326 => to_slv(opcode_type, 16#10#),
      327 => to_slv(opcode_type, 16#0C#),
      328 => to_slv(opcode_type, 16#06#),
      329 => to_slv(opcode_type, 16#09#),
      330 => to_slv(opcode_type, 16#0A#),
      331 => to_slv(opcode_type, 16#0C#),
      332 => to_slv(opcode_type, 16#08#),
      333 => to_slv(opcode_type, 16#0C#),
      334 => to_slv(opcode_type, 16#0B#),
      335 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#07#),
      353 => to_slv(opcode_type, 16#05#),
      354 => to_slv(opcode_type, 16#07#),
      355 => to_slv(opcode_type, 16#04#),
      356 => to_slv(opcode_type, 16#10#),
      357 => to_slv(opcode_type, 16#05#),
      358 => to_slv(opcode_type, 16#11#),
      359 => to_slv(opcode_type, 16#06#),
      360 => to_slv(opcode_type, 16#06#),
      361 => to_slv(opcode_type, 16#07#),
      362 => to_slv(opcode_type, 16#0A#),
      363 => to_slv(opcode_type, 16#10#),
      364 => to_slv(opcode_type, 16#04#),
      365 => to_slv(opcode_type, 16#D2#),
      366 => to_slv(opcode_type, 16#9A#),
      367 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#01#),
      385 => to_slv(opcode_type, 16#08#),
      386 => to_slv(opcode_type, 16#09#),
      387 => to_slv(opcode_type, 16#04#),
      388 => to_slv(opcode_type, 16#0B#),
      389 => to_slv(opcode_type, 16#06#),
      390 => to_slv(opcode_type, 16#11#),
      391 => to_slv(opcode_type, 16#25#),
      392 => to_slv(opcode_type, 16#09#),
      393 => to_slv(opcode_type, 16#07#),
      394 => to_slv(opcode_type, 16#11#),
      395 => to_slv(opcode_type, 16#0A#),
      396 => to_slv(opcode_type, 16#09#),
      397 => to_slv(opcode_type, 16#11#),
      398 => to_slv(opcode_type, 16#10#),
      399 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#07#),
      417 => to_slv(opcode_type, 16#03#),
      418 => to_slv(opcode_type, 16#04#),
      419 => to_slv(opcode_type, 16#02#),
      420 => to_slv(opcode_type, 16#11#),
      421 => to_slv(opcode_type, 16#06#),
      422 => to_slv(opcode_type, 16#07#),
      423 => to_slv(opcode_type, 16#07#),
      424 => to_slv(opcode_type, 16#10#),
      425 => to_slv(opcode_type, 16#10#),
      426 => to_slv(opcode_type, 16#03#),
      427 => to_slv(opcode_type, 16#C1#),
      428 => to_slv(opcode_type, 16#02#),
      429 => to_slv(opcode_type, 16#02#),
      430 => to_slv(opcode_type, 16#0B#),
      431 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#04#),
      449 => to_slv(opcode_type, 16#06#),
      450 => to_slv(opcode_type, 16#07#),
      451 => to_slv(opcode_type, 16#01#),
      452 => to_slv(opcode_type, 16#27#),
      453 => to_slv(opcode_type, 16#09#),
      454 => to_slv(opcode_type, 16#0F#),
      455 => to_slv(opcode_type, 16#10#),
      456 => to_slv(opcode_type, 16#08#),
      457 => to_slv(opcode_type, 16#06#),
      458 => to_slv(opcode_type, 16#0C#),
      459 => to_slv(opcode_type, 16#10#),
      460 => to_slv(opcode_type, 16#07#),
      461 => to_slv(opcode_type, 16#0A#),
      462 => to_slv(opcode_type, 16#0E#),
      463 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#06#),
      481 => to_slv(opcode_type, 16#06#),
      482 => to_slv(opcode_type, 16#01#),
      483 => to_slv(opcode_type, 16#09#),
      484 => to_slv(opcode_type, 16#89#),
      485 => to_slv(opcode_type, 16#0E#),
      486 => to_slv(opcode_type, 16#01#),
      487 => to_slv(opcode_type, 16#09#),
      488 => to_slv(opcode_type, 16#0B#),
      489 => to_slv(opcode_type, 16#0C#),
      490 => to_slv(opcode_type, 16#08#),
      491 => to_slv(opcode_type, 16#06#),
      492 => to_slv(opcode_type, 16#0F#),
      493 => to_slv(opcode_type, 16#0A#),
      494 => to_slv(opcode_type, 16#0A#),
      495 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#07#),
      513 => to_slv(opcode_type, 16#02#),
      514 => to_slv(opcode_type, 16#08#),
      515 => to_slv(opcode_type, 16#03#),
      516 => to_slv(opcode_type, 16#0A#),
      517 => to_slv(opcode_type, 16#03#),
      518 => to_slv(opcode_type, 16#0F#),
      519 => to_slv(opcode_type, 16#08#),
      520 => to_slv(opcode_type, 16#08#),
      521 => to_slv(opcode_type, 16#01#),
      522 => to_slv(opcode_type, 16#11#),
      523 => to_slv(opcode_type, 16#01#),
      524 => to_slv(opcode_type, 16#B4#),
      525 => to_slv(opcode_type, 16#03#),
      526 => to_slv(opcode_type, 16#11#),
      527 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#04#),
      545 => to_slv(opcode_type, 16#08#),
      546 => to_slv(opcode_type, 16#08#),
      547 => to_slv(opcode_type, 16#04#),
      548 => to_slv(opcode_type, 16#0C#),
      549 => to_slv(opcode_type, 16#08#),
      550 => to_slv(opcode_type, 16#0D#),
      551 => to_slv(opcode_type, 16#11#),
      552 => to_slv(opcode_type, 16#09#),
      553 => to_slv(opcode_type, 16#06#),
      554 => to_slv(opcode_type, 16#11#),
      555 => to_slv(opcode_type, 16#0B#),
      556 => to_slv(opcode_type, 16#08#),
      557 => to_slv(opcode_type, 16#0A#),
      558 => to_slv(opcode_type, 16#10#),
      559 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#06#),
      577 => to_slv(opcode_type, 16#01#),
      578 => to_slv(opcode_type, 16#06#),
      579 => to_slv(opcode_type, 16#08#),
      580 => to_slv(opcode_type, 16#0D#),
      581 => to_slv(opcode_type, 16#0D#),
      582 => to_slv(opcode_type, 16#05#),
      583 => to_slv(opcode_type, 16#0E#),
      584 => to_slv(opcode_type, 16#04#),
      585 => to_slv(opcode_type, 16#08#),
      586 => to_slv(opcode_type, 16#06#),
      587 => to_slv(opcode_type, 16#D4#),
      588 => to_slv(opcode_type, 16#10#),
      589 => to_slv(opcode_type, 16#02#),
      590 => to_slv(opcode_type, 16#93#),
      591 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#06#),
      609 => to_slv(opcode_type, 16#06#),
      610 => to_slv(opcode_type, 16#07#),
      611 => to_slv(opcode_type, 16#08#),
      612 => to_slv(opcode_type, 16#11#),
      613 => to_slv(opcode_type, 16#0F#),
      614 => to_slv(opcode_type, 16#09#),
      615 => to_slv(opcode_type, 16#10#),
      616 => to_slv(opcode_type, 16#0C#),
      617 => to_slv(opcode_type, 16#07#),
      618 => to_slv(opcode_type, 16#08#),
      619 => to_slv(opcode_type, 16#0F#),
      620 => to_slv(opcode_type, 16#0F#),
      621 => to_slv(opcode_type, 16#0E#),
      622 => to_slv(opcode_type, 16#0A#),
      623 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#09#),
      641 => to_slv(opcode_type, 16#07#),
      642 => to_slv(opcode_type, 16#09#),
      643 => to_slv(opcode_type, 16#04#),
      644 => to_slv(opcode_type, 16#0D#),
      645 => to_slv(opcode_type, 16#06#),
      646 => to_slv(opcode_type, 16#10#),
      647 => to_slv(opcode_type, 16#0C#),
      648 => to_slv(opcode_type, 16#05#),
      649 => to_slv(opcode_type, 16#08#),
      650 => to_slv(opcode_type, 16#11#),
      651 => to_slv(opcode_type, 16#10#),
      652 => to_slv(opcode_type, 16#02#),
      653 => to_slv(opcode_type, 16#01#),
      654 => to_slv(opcode_type, 16#0C#),
      655 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#04#),
      673 => to_slv(opcode_type, 16#09#),
      674 => to_slv(opcode_type, 16#08#),
      675 => to_slv(opcode_type, 16#02#),
      676 => to_slv(opcode_type, 16#0A#),
      677 => to_slv(opcode_type, 16#07#),
      678 => to_slv(opcode_type, 16#0A#),
      679 => to_slv(opcode_type, 16#0E#),
      680 => to_slv(opcode_type, 16#09#),
      681 => to_slv(opcode_type, 16#07#),
      682 => to_slv(opcode_type, 16#0D#),
      683 => to_slv(opcode_type, 16#0E#),
      684 => to_slv(opcode_type, 16#07#),
      685 => to_slv(opcode_type, 16#0B#),
      686 => to_slv(opcode_type, 16#0D#),
      687 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#04#),
      705 => to_slv(opcode_type, 16#09#),
      706 => to_slv(opcode_type, 16#08#),
      707 => to_slv(opcode_type, 16#07#),
      708 => to_slv(opcode_type, 16#6D#),
      709 => to_slv(opcode_type, 16#0D#),
      710 => to_slv(opcode_type, 16#02#),
      711 => to_slv(opcode_type, 16#0D#),
      712 => to_slv(opcode_type, 16#06#),
      713 => to_slv(opcode_type, 16#09#),
      714 => to_slv(opcode_type, 16#0D#),
      715 => to_slv(opcode_type, 16#10#),
      716 => to_slv(opcode_type, 16#07#),
      717 => to_slv(opcode_type, 16#10#),
      718 => to_slv(opcode_type, 16#0B#),
      719 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#02#),
      737 => to_slv(opcode_type, 16#09#),
      738 => to_slv(opcode_type, 16#08#),
      739 => to_slv(opcode_type, 16#06#),
      740 => to_slv(opcode_type, 16#0C#),
      741 => to_slv(opcode_type, 16#11#),
      742 => to_slv(opcode_type, 16#04#),
      743 => to_slv(opcode_type, 16#0A#),
      744 => to_slv(opcode_type, 16#08#),
      745 => to_slv(opcode_type, 16#08#),
      746 => to_slv(opcode_type, 16#0E#),
      747 => to_slv(opcode_type, 16#11#),
      748 => to_slv(opcode_type, 16#06#),
      749 => to_slv(opcode_type, 16#0A#),
      750 => to_slv(opcode_type, 16#0B#),
      751 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#01#),
      769 => to_slv(opcode_type, 16#07#),
      770 => to_slv(opcode_type, 16#07#),
      771 => to_slv(opcode_type, 16#04#),
      772 => to_slv(opcode_type, 16#10#),
      773 => to_slv(opcode_type, 16#08#),
      774 => to_slv(opcode_type, 16#0B#),
      775 => to_slv(opcode_type, 16#0E#),
      776 => to_slv(opcode_type, 16#08#),
      777 => to_slv(opcode_type, 16#07#),
      778 => to_slv(opcode_type, 16#0C#),
      779 => to_slv(opcode_type, 16#0B#),
      780 => to_slv(opcode_type, 16#07#),
      781 => to_slv(opcode_type, 16#0D#),
      782 => to_slv(opcode_type, 16#0F#),
      783 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#08#),
      801 => to_slv(opcode_type, 16#02#),
      802 => to_slv(opcode_type, 16#09#),
      803 => to_slv(opcode_type, 16#05#),
      804 => to_slv(opcode_type, 16#0E#),
      805 => to_slv(opcode_type, 16#03#),
      806 => to_slv(opcode_type, 16#0B#),
      807 => to_slv(opcode_type, 16#01#),
      808 => to_slv(opcode_type, 16#09#),
      809 => to_slv(opcode_type, 16#09#),
      810 => to_slv(opcode_type, 16#0F#),
      811 => to_slv(opcode_type, 16#10#),
      812 => to_slv(opcode_type, 16#08#),
      813 => to_slv(opcode_type, 16#0B#),
      814 => to_slv(opcode_type, 16#0F#),
      815 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#04#),
      833 => to_slv(opcode_type, 16#07#),
      834 => to_slv(opcode_type, 16#06#),
      835 => to_slv(opcode_type, 16#06#),
      836 => to_slv(opcode_type, 16#0A#),
      837 => to_slv(opcode_type, 16#0C#),
      838 => to_slv(opcode_type, 16#06#),
      839 => to_slv(opcode_type, 16#0B#),
      840 => to_slv(opcode_type, 16#13#),
      841 => to_slv(opcode_type, 16#06#),
      842 => to_slv(opcode_type, 16#05#),
      843 => to_slv(opcode_type, 16#0F#),
      844 => to_slv(opcode_type, 16#06#),
      845 => to_slv(opcode_type, 16#0F#),
      846 => to_slv(opcode_type, 16#0E#),
      847 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#07#),
      865 => to_slv(opcode_type, 16#05#),
      866 => to_slv(opcode_type, 16#06#),
      867 => to_slv(opcode_type, 16#04#),
      868 => to_slv(opcode_type, 16#0B#),
      869 => to_slv(opcode_type, 16#04#),
      870 => to_slv(opcode_type, 16#0D#),
      871 => to_slv(opcode_type, 16#09#),
      872 => to_slv(opcode_type, 16#08#),
      873 => to_slv(opcode_type, 16#04#),
      874 => to_slv(opcode_type, 16#8B#),
      875 => to_slv(opcode_type, 16#06#),
      876 => to_slv(opcode_type, 16#BC#),
      877 => to_slv(opcode_type, 16#0B#),
      878 => to_slv(opcode_type, 16#0C#),
      879 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#09#),
      898 => to_slv(opcode_type, 16#02#),
      899 => to_slv(opcode_type, 16#04#),
      900 => to_slv(opcode_type, 16#D9#),
      901 => to_slv(opcode_type, 16#03#),
      902 => to_slv(opcode_type, 16#07#),
      903 => to_slv(opcode_type, 16#0A#),
      904 => to_slv(opcode_type, 16#0A#),
      905 => to_slv(opcode_type, 16#06#),
      906 => to_slv(opcode_type, 16#06#),
      907 => to_slv(opcode_type, 16#05#),
      908 => to_slv(opcode_type, 16#0C#),
      909 => to_slv(opcode_type, 16#11#),
      910 => to_slv(opcode_type, 16#10#),
      911 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#04#),
      929 => to_slv(opcode_type, 16#08#),
      930 => to_slv(opcode_type, 16#08#),
      931 => to_slv(opcode_type, 16#08#),
      932 => to_slv(opcode_type, 16#E0#),
      933 => to_slv(opcode_type, 16#0F#),
      934 => to_slv(opcode_type, 16#07#),
      935 => to_slv(opcode_type, 16#0B#),
      936 => to_slv(opcode_type, 16#10#),
      937 => to_slv(opcode_type, 16#06#),
      938 => to_slv(opcode_type, 16#04#),
      939 => to_slv(opcode_type, 16#0F#),
      940 => to_slv(opcode_type, 16#07#),
      941 => to_slv(opcode_type, 16#0B#),
      942 => to_slv(opcode_type, 16#0A#),
      943 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#05#),
      962 => to_slv(opcode_type, 16#02#),
      963 => to_slv(opcode_type, 16#04#),
      964 => to_slv(opcode_type, 16#0F#),
      965 => to_slv(opcode_type, 16#06#),
      966 => to_slv(opcode_type, 16#09#),
      967 => to_slv(opcode_type, 16#02#),
      968 => to_slv(opcode_type, 16#D2#),
      969 => to_slv(opcode_type, 16#02#),
      970 => to_slv(opcode_type, 16#0D#),
      971 => to_slv(opcode_type, 16#09#),
      972 => to_slv(opcode_type, 16#05#),
      973 => to_slv(opcode_type, 16#0E#),
      974 => to_slv(opcode_type, 16#19#),
      975 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#08#),
      993 => to_slv(opcode_type, 16#03#),
      994 => to_slv(opcode_type, 16#09#),
      995 => to_slv(opcode_type, 16#01#),
      996 => to_slv(opcode_type, 16#C5#),
      997 => to_slv(opcode_type, 16#04#),
      998 => to_slv(opcode_type, 16#0B#),
      999 => to_slv(opcode_type, 16#03#),
      1000 => to_slv(opcode_type, 16#08#),
      1001 => to_slv(opcode_type, 16#09#),
      1002 => to_slv(opcode_type, 16#10#),
      1003 => to_slv(opcode_type, 16#11#),
      1004 => to_slv(opcode_type, 16#06#),
      1005 => to_slv(opcode_type, 16#0B#),
      1006 => to_slv(opcode_type, 16#0E#),
      1007 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#07#),
      1025 => to_slv(opcode_type, 16#08#),
      1026 => to_slv(opcode_type, 16#02#),
      1027 => to_slv(opcode_type, 16#03#),
      1028 => to_slv(opcode_type, 16#6F#),
      1029 => to_slv(opcode_type, 16#05#),
      1030 => to_slv(opcode_type, 16#05#),
      1031 => to_slv(opcode_type, 16#0D#),
      1032 => to_slv(opcode_type, 16#06#),
      1033 => to_slv(opcode_type, 16#04#),
      1034 => to_slv(opcode_type, 16#02#),
      1035 => to_slv(opcode_type, 16#0E#),
      1036 => to_slv(opcode_type, 16#03#),
      1037 => to_slv(opcode_type, 16#01#),
      1038 => to_slv(opcode_type, 16#0F#),
      1039 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#02#),
      1057 => to_slv(opcode_type, 16#06#),
      1058 => to_slv(opcode_type, 16#09#),
      1059 => to_slv(opcode_type, 16#06#),
      1060 => to_slv(opcode_type, 16#0A#),
      1061 => to_slv(opcode_type, 16#0A#),
      1062 => to_slv(opcode_type, 16#04#),
      1063 => to_slv(opcode_type, 16#0A#),
      1064 => to_slv(opcode_type, 16#08#),
      1065 => to_slv(opcode_type, 16#09#),
      1066 => to_slv(opcode_type, 16#0B#),
      1067 => to_slv(opcode_type, 16#0B#),
      1068 => to_slv(opcode_type, 16#07#),
      1069 => to_slv(opcode_type, 16#0B#),
      1070 => to_slv(opcode_type, 16#10#),
      1071 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#03#),
      1089 => to_slv(opcode_type, 16#07#),
      1090 => to_slv(opcode_type, 16#08#),
      1091 => to_slv(opcode_type, 16#08#),
      1092 => to_slv(opcode_type, 16#0F#),
      1093 => to_slv(opcode_type, 16#D0#),
      1094 => to_slv(opcode_type, 16#07#),
      1095 => to_slv(opcode_type, 16#11#),
      1096 => to_slv(opcode_type, 16#10#),
      1097 => to_slv(opcode_type, 16#09#),
      1098 => to_slv(opcode_type, 16#05#),
      1099 => to_slv(opcode_type, 16#11#),
      1100 => to_slv(opcode_type, 16#08#),
      1101 => to_slv(opcode_type, 16#11#),
      1102 => to_slv(opcode_type, 16#10#),
      1103 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#05#),
      1121 => to_slv(opcode_type, 16#08#),
      1122 => to_slv(opcode_type, 16#06#),
      1123 => to_slv(opcode_type, 16#01#),
      1124 => to_slv(opcode_type, 16#0F#),
      1125 => to_slv(opcode_type, 16#08#),
      1126 => to_slv(opcode_type, 16#C0#),
      1127 => to_slv(opcode_type, 16#0C#),
      1128 => to_slv(opcode_type, 16#09#),
      1129 => to_slv(opcode_type, 16#06#),
      1130 => to_slv(opcode_type, 16#11#),
      1131 => to_slv(opcode_type, 16#E4#),
      1132 => to_slv(opcode_type, 16#09#),
      1133 => to_slv(opcode_type, 16#0D#),
      1134 => to_slv(opcode_type, 16#0F#),
      1135 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#04#),
      1153 => to_slv(opcode_type, 16#07#),
      1154 => to_slv(opcode_type, 16#07#),
      1155 => to_slv(opcode_type, 16#05#),
      1156 => to_slv(opcode_type, 16#0C#),
      1157 => to_slv(opcode_type, 16#07#),
      1158 => to_slv(opcode_type, 16#10#),
      1159 => to_slv(opcode_type, 16#0B#),
      1160 => to_slv(opcode_type, 16#08#),
      1161 => to_slv(opcode_type, 16#07#),
      1162 => to_slv(opcode_type, 16#0A#),
      1163 => to_slv(opcode_type, 16#0E#),
      1164 => to_slv(opcode_type, 16#07#),
      1165 => to_slv(opcode_type, 16#11#),
      1166 => to_slv(opcode_type, 16#0D#),
      1167 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#09#),
      1185 => to_slv(opcode_type, 16#03#),
      1186 => to_slv(opcode_type, 16#03#),
      1187 => to_slv(opcode_type, 16#03#),
      1188 => to_slv(opcode_type, 16#11#),
      1189 => to_slv(opcode_type, 16#06#),
      1190 => to_slv(opcode_type, 16#03#),
      1191 => to_slv(opcode_type, 16#06#),
      1192 => to_slv(opcode_type, 16#0C#),
      1193 => to_slv(opcode_type, 16#10#),
      1194 => to_slv(opcode_type, 16#08#),
      1195 => to_slv(opcode_type, 16#03#),
      1196 => to_slv(opcode_type, 16#0C#),
      1197 => to_slv(opcode_type, 16#03#),
      1198 => to_slv(opcode_type, 16#0F#),
      1199 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#08#),
      1217 => to_slv(opcode_type, 16#01#),
      1218 => to_slv(opcode_type, 16#07#),
      1219 => to_slv(opcode_type, 16#01#),
      1220 => to_slv(opcode_type, 16#0E#),
      1221 => to_slv(opcode_type, 16#05#),
      1222 => to_slv(opcode_type, 16#0C#),
      1223 => to_slv(opcode_type, 16#01#),
      1224 => to_slv(opcode_type, 16#09#),
      1225 => to_slv(opcode_type, 16#08#),
      1226 => to_slv(opcode_type, 16#11#),
      1227 => to_slv(opcode_type, 16#0A#),
      1228 => to_slv(opcode_type, 16#07#),
      1229 => to_slv(opcode_type, 16#AD#),
      1230 => to_slv(opcode_type, 16#0B#),
      1231 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#03#),
      1249 => to_slv(opcode_type, 16#09#),
      1250 => to_slv(opcode_type, 16#08#),
      1251 => to_slv(opcode_type, 16#09#),
      1252 => to_slv(opcode_type, 16#11#),
      1253 => to_slv(opcode_type, 16#0A#),
      1254 => to_slv(opcode_type, 16#04#),
      1255 => to_slv(opcode_type, 16#0A#),
      1256 => to_slv(opcode_type, 16#06#),
      1257 => to_slv(opcode_type, 16#08#),
      1258 => to_slv(opcode_type, 16#11#),
      1259 => to_slv(opcode_type, 16#0C#),
      1260 => to_slv(opcode_type, 16#07#),
      1261 => to_slv(opcode_type, 16#0F#),
      1262 => to_slv(opcode_type, 16#0E#),
      1263 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#07#),
      1281 => to_slv(opcode_type, 16#01#),
      1282 => to_slv(opcode_type, 16#09#),
      1283 => to_slv(opcode_type, 16#09#),
      1284 => to_slv(opcode_type, 16#0E#),
      1285 => to_slv(opcode_type, 16#0A#),
      1286 => to_slv(opcode_type, 16#09#),
      1287 => to_slv(opcode_type, 16#C5#),
      1288 => to_slv(opcode_type, 16#58#),
      1289 => to_slv(opcode_type, 16#08#),
      1290 => to_slv(opcode_type, 16#04#),
      1291 => to_slv(opcode_type, 16#02#),
      1292 => to_slv(opcode_type, 16#0D#),
      1293 => to_slv(opcode_type, 16#02#),
      1294 => to_slv(opcode_type, 16#0E#),
      1295 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#06#),
      1313 => to_slv(opcode_type, 16#04#),
      1314 => to_slv(opcode_type, 16#05#),
      1315 => to_slv(opcode_type, 16#09#),
      1316 => to_slv(opcode_type, 16#0A#),
      1317 => to_slv(opcode_type, 16#0C#),
      1318 => to_slv(opcode_type, 16#06#),
      1319 => to_slv(opcode_type, 16#01#),
      1320 => to_slv(opcode_type, 16#06#),
      1321 => to_slv(opcode_type, 16#11#),
      1322 => to_slv(opcode_type, 16#0D#),
      1323 => to_slv(opcode_type, 16#01#),
      1324 => to_slv(opcode_type, 16#07#),
      1325 => to_slv(opcode_type, 16#10#),
      1326 => to_slv(opcode_type, 16#0A#),
      1327 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#09#),
      1345 => to_slv(opcode_type, 16#02#),
      1346 => to_slv(opcode_type, 16#07#),
      1347 => to_slv(opcode_type, 16#09#),
      1348 => to_slv(opcode_type, 16#B0#),
      1349 => to_slv(opcode_type, 16#0D#),
      1350 => to_slv(opcode_type, 16#07#),
      1351 => to_slv(opcode_type, 16#6D#),
      1352 => to_slv(opcode_type, 16#ED#),
      1353 => to_slv(opcode_type, 16#08#),
      1354 => to_slv(opcode_type, 16#05#),
      1355 => to_slv(opcode_type, 16#05#),
      1356 => to_slv(opcode_type, 16#0D#),
      1357 => to_slv(opcode_type, 16#05#),
      1358 => to_slv(opcode_type, 16#11#),
      1359 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#02#),
      1377 => to_slv(opcode_type, 16#08#),
      1378 => to_slv(opcode_type, 16#08#),
      1379 => to_slv(opcode_type, 16#03#),
      1380 => to_slv(opcode_type, 16#0F#),
      1381 => to_slv(opcode_type, 16#06#),
      1382 => to_slv(opcode_type, 16#0B#),
      1383 => to_slv(opcode_type, 16#0B#),
      1384 => to_slv(opcode_type, 16#09#),
      1385 => to_slv(opcode_type, 16#08#),
      1386 => to_slv(opcode_type, 16#0E#),
      1387 => to_slv(opcode_type, 16#C3#),
      1388 => to_slv(opcode_type, 16#06#),
      1389 => to_slv(opcode_type, 16#0B#),
      1390 => to_slv(opcode_type, 16#0B#),
      1391 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#04#),
      1409 => to_slv(opcode_type, 16#06#),
      1410 => to_slv(opcode_type, 16#09#),
      1411 => to_slv(opcode_type, 16#01#),
      1412 => to_slv(opcode_type, 16#F7#),
      1413 => to_slv(opcode_type, 16#06#),
      1414 => to_slv(opcode_type, 16#0B#),
      1415 => to_slv(opcode_type, 16#0A#),
      1416 => to_slv(opcode_type, 16#09#),
      1417 => to_slv(opcode_type, 16#06#),
      1418 => to_slv(opcode_type, 16#10#),
      1419 => to_slv(opcode_type, 16#0F#),
      1420 => to_slv(opcode_type, 16#06#),
      1421 => to_slv(opcode_type, 16#11#),
      1422 => to_slv(opcode_type, 16#0D#),
      1423 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#02#),
      1441 => to_slv(opcode_type, 16#09#),
      1442 => to_slv(opcode_type, 16#07#),
      1443 => to_slv(opcode_type, 16#07#),
      1444 => to_slv(opcode_type, 16#0C#),
      1445 => to_slv(opcode_type, 16#13#),
      1446 => to_slv(opcode_type, 16#04#),
      1447 => to_slv(opcode_type, 16#0F#),
      1448 => to_slv(opcode_type, 16#09#),
      1449 => to_slv(opcode_type, 16#07#),
      1450 => to_slv(opcode_type, 16#5B#),
      1451 => to_slv(opcode_type, 16#0F#),
      1452 => to_slv(opcode_type, 16#09#),
      1453 => to_slv(opcode_type, 16#0A#),
      1454 => to_slv(opcode_type, 16#11#),
      1455 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#07#),
      1473 => to_slv(opcode_type, 16#09#),
      1474 => to_slv(opcode_type, 16#05#),
      1475 => to_slv(opcode_type, 16#08#),
      1476 => to_slv(opcode_type, 16#10#),
      1477 => to_slv(opcode_type, 16#0B#),
      1478 => to_slv(opcode_type, 16#06#),
      1479 => to_slv(opcode_type, 16#07#),
      1480 => to_slv(opcode_type, 16#2C#),
      1481 => to_slv(opcode_type, 16#10#),
      1482 => to_slv(opcode_type, 16#08#),
      1483 => to_slv(opcode_type, 16#0D#),
      1484 => to_slv(opcode_type, 16#10#),
      1485 => to_slv(opcode_type, 16#04#),
      1486 => to_slv(opcode_type, 16#0B#),
      1487 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#04#),
      1505 => to_slv(opcode_type, 16#08#),
      1506 => to_slv(opcode_type, 16#09#),
      1507 => to_slv(opcode_type, 16#01#),
      1508 => to_slv(opcode_type, 16#10#),
      1509 => to_slv(opcode_type, 16#06#),
      1510 => to_slv(opcode_type, 16#0F#),
      1511 => to_slv(opcode_type, 16#0C#),
      1512 => to_slv(opcode_type, 16#08#),
      1513 => to_slv(opcode_type, 16#07#),
      1514 => to_slv(opcode_type, 16#11#),
      1515 => to_slv(opcode_type, 16#10#),
      1516 => to_slv(opcode_type, 16#08#),
      1517 => to_slv(opcode_type, 16#0A#),
      1518 => to_slv(opcode_type, 16#10#),
      1519 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#05#),
      1537 => to_slv(opcode_type, 16#09#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#09#),
      1540 => to_slv(opcode_type, 16#0D#),
      1541 => to_slv(opcode_type, 16#9A#),
      1542 => to_slv(opcode_type, 16#02#),
      1543 => to_slv(opcode_type, 16#0B#),
      1544 => to_slv(opcode_type, 16#07#),
      1545 => to_slv(opcode_type, 16#06#),
      1546 => to_slv(opcode_type, 16#0E#),
      1547 => to_slv(opcode_type, 16#11#),
      1548 => to_slv(opcode_type, 16#07#),
      1549 => to_slv(opcode_type, 16#0C#),
      1550 => to_slv(opcode_type, 16#0A#),
      1551 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#06#),
      1569 => to_slv(opcode_type, 16#03#),
      1570 => to_slv(opcode_type, 16#03#),
      1571 => to_slv(opcode_type, 16#07#),
      1572 => to_slv(opcode_type, 16#0D#),
      1573 => to_slv(opcode_type, 16#10#),
      1574 => to_slv(opcode_type, 16#06#),
      1575 => to_slv(opcode_type, 16#07#),
      1576 => to_slv(opcode_type, 16#05#),
      1577 => to_slv(opcode_type, 16#0C#),
      1578 => to_slv(opcode_type, 16#08#),
      1579 => to_slv(opcode_type, 16#11#),
      1580 => to_slv(opcode_type, 16#0E#),
      1581 => to_slv(opcode_type, 16#04#),
      1582 => to_slv(opcode_type, 16#11#),
      1583 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#07#),
      1601 => to_slv(opcode_type, 16#01#),
      1602 => to_slv(opcode_type, 16#08#),
      1603 => to_slv(opcode_type, 16#03#),
      1604 => to_slv(opcode_type, 16#0F#),
      1605 => to_slv(opcode_type, 16#05#),
      1606 => to_slv(opcode_type, 16#10#),
      1607 => to_slv(opcode_type, 16#01#),
      1608 => to_slv(opcode_type, 16#09#),
      1609 => to_slv(opcode_type, 16#09#),
      1610 => to_slv(opcode_type, 16#0C#),
      1611 => to_slv(opcode_type, 16#0D#),
      1612 => to_slv(opcode_type, 16#08#),
      1613 => to_slv(opcode_type, 16#0D#),
      1614 => to_slv(opcode_type, 16#0C#),
      1615 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#01#),
      1633 => to_slv(opcode_type, 16#07#),
      1634 => to_slv(opcode_type, 16#08#),
      1635 => to_slv(opcode_type, 16#05#),
      1636 => to_slv(opcode_type, 16#0A#),
      1637 => to_slv(opcode_type, 16#08#),
      1638 => to_slv(opcode_type, 16#0C#),
      1639 => to_slv(opcode_type, 16#0A#),
      1640 => to_slv(opcode_type, 16#06#),
      1641 => to_slv(opcode_type, 16#09#),
      1642 => to_slv(opcode_type, 16#0A#),
      1643 => to_slv(opcode_type, 16#0F#),
      1644 => to_slv(opcode_type, 16#08#),
      1645 => to_slv(opcode_type, 16#10#),
      1646 => to_slv(opcode_type, 16#0B#),
      1647 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#06#),
      1665 => to_slv(opcode_type, 16#04#),
      1666 => to_slv(opcode_type, 16#06#),
      1667 => to_slv(opcode_type, 16#01#),
      1668 => to_slv(opcode_type, 16#11#),
      1669 => to_slv(opcode_type, 16#01#),
      1670 => to_slv(opcode_type, 16#0B#),
      1671 => to_slv(opcode_type, 16#06#),
      1672 => to_slv(opcode_type, 16#09#),
      1673 => to_slv(opcode_type, 16#03#),
      1674 => to_slv(opcode_type, 16#0A#),
      1675 => to_slv(opcode_type, 16#06#),
      1676 => to_slv(opcode_type, 16#10#),
      1677 => to_slv(opcode_type, 16#11#),
      1678 => to_slv(opcode_type, 16#81#),
      1679 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#09#),
      1697 => to_slv(opcode_type, 16#01#),
      1698 => to_slv(opcode_type, 16#05#),
      1699 => to_slv(opcode_type, 16#01#),
      1700 => to_slv(opcode_type, 16#0D#),
      1701 => to_slv(opcode_type, 16#09#),
      1702 => to_slv(opcode_type, 16#04#),
      1703 => to_slv(opcode_type, 16#02#),
      1704 => to_slv(opcode_type, 16#0C#),
      1705 => to_slv(opcode_type, 16#07#),
      1706 => to_slv(opcode_type, 16#06#),
      1707 => to_slv(opcode_type, 16#0D#),
      1708 => to_slv(opcode_type, 16#0F#),
      1709 => to_slv(opcode_type, 16#04#),
      1710 => to_slv(opcode_type, 16#0A#),
      1711 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#05#),
      1729 => to_slv(opcode_type, 16#08#),
      1730 => to_slv(opcode_type, 16#07#),
      1731 => to_slv(opcode_type, 16#01#),
      1732 => to_slv(opcode_type, 16#0B#),
      1733 => to_slv(opcode_type, 16#09#),
      1734 => to_slv(opcode_type, 16#CC#),
      1735 => to_slv(opcode_type, 16#10#),
      1736 => to_slv(opcode_type, 16#09#),
      1737 => to_slv(opcode_type, 16#06#),
      1738 => to_slv(opcode_type, 16#0C#),
      1739 => to_slv(opcode_type, 16#0A#),
      1740 => to_slv(opcode_type, 16#06#),
      1741 => to_slv(opcode_type, 16#0E#),
      1742 => to_slv(opcode_type, 16#0D#),
      1743 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#07#),
      1761 => to_slv(opcode_type, 16#09#),
      1762 => to_slv(opcode_type, 16#05#),
      1763 => to_slv(opcode_type, 16#07#),
      1764 => to_slv(opcode_type, 16#0B#),
      1765 => to_slv(opcode_type, 16#0F#),
      1766 => to_slv(opcode_type, 16#09#),
      1767 => to_slv(opcode_type, 16#07#),
      1768 => to_slv(opcode_type, 16#0D#),
      1769 => to_slv(opcode_type, 16#0D#),
      1770 => to_slv(opcode_type, 16#02#),
      1771 => to_slv(opcode_type, 16#0E#),
      1772 => to_slv(opcode_type, 16#05#),
      1773 => to_slv(opcode_type, 16#01#),
      1774 => to_slv(opcode_type, 16#0E#),
      1775 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#06#),
      1793 => to_slv(opcode_type, 16#06#),
      1794 => to_slv(opcode_type, 16#04#),
      1795 => to_slv(opcode_type, 16#02#),
      1796 => to_slv(opcode_type, 16#0B#),
      1797 => to_slv(opcode_type, 16#02#),
      1798 => to_slv(opcode_type, 16#09#),
      1799 => to_slv(opcode_type, 16#0A#),
      1800 => to_slv(opcode_type, 16#0A#),
      1801 => to_slv(opcode_type, 16#01#),
      1802 => to_slv(opcode_type, 16#06#),
      1803 => to_slv(opcode_type, 16#07#),
      1804 => to_slv(opcode_type, 16#0D#),
      1805 => to_slv(opcode_type, 16#11#),
      1806 => to_slv(opcode_type, 16#0A#),
      1807 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#01#),
      1825 => to_slv(opcode_type, 16#08#),
      1826 => to_slv(opcode_type, 16#06#),
      1827 => to_slv(opcode_type, 16#02#),
      1828 => to_slv(opcode_type, 16#0B#),
      1829 => to_slv(opcode_type, 16#09#),
      1830 => to_slv(opcode_type, 16#0E#),
      1831 => to_slv(opcode_type, 16#11#),
      1832 => to_slv(opcode_type, 16#08#),
      1833 => to_slv(opcode_type, 16#08#),
      1834 => to_slv(opcode_type, 16#0C#),
      1835 => to_slv(opcode_type, 16#95#),
      1836 => to_slv(opcode_type, 16#06#),
      1837 => to_slv(opcode_type, 16#10#),
      1838 => to_slv(opcode_type, 16#0B#),
      1839 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#06#),
      1857 => to_slv(opcode_type, 16#04#),
      1858 => to_slv(opcode_type, 16#01#),
      1859 => to_slv(opcode_type, 16#06#),
      1860 => to_slv(opcode_type, 16#0B#),
      1861 => to_slv(opcode_type, 16#11#),
      1862 => to_slv(opcode_type, 16#09#),
      1863 => to_slv(opcode_type, 16#04#),
      1864 => to_slv(opcode_type, 16#03#),
      1865 => to_slv(opcode_type, 16#11#),
      1866 => to_slv(opcode_type, 16#07#),
      1867 => to_slv(opcode_type, 16#09#),
      1868 => to_slv(opcode_type, 16#C2#),
      1869 => to_slv(opcode_type, 16#0C#),
      1870 => to_slv(opcode_type, 16#0F#),
      1871 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#02#),
      1889 => to_slv(opcode_type, 16#09#),
      1890 => to_slv(opcode_type, 16#06#),
      1891 => to_slv(opcode_type, 16#01#),
      1892 => to_slv(opcode_type, 16#0E#),
      1893 => to_slv(opcode_type, 16#08#),
      1894 => to_slv(opcode_type, 16#0A#),
      1895 => to_slv(opcode_type, 16#0E#),
      1896 => to_slv(opcode_type, 16#09#),
      1897 => to_slv(opcode_type, 16#08#),
      1898 => to_slv(opcode_type, 16#0C#),
      1899 => to_slv(opcode_type, 16#0C#),
      1900 => to_slv(opcode_type, 16#09#),
      1901 => to_slv(opcode_type, 16#0B#),
      1902 => to_slv(opcode_type, 16#0E#),
      1903 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#04#),
      1921 => to_slv(opcode_type, 16#08#),
      1922 => to_slv(opcode_type, 16#09#),
      1923 => to_slv(opcode_type, 16#07#),
      1924 => to_slv(opcode_type, 16#10#),
      1925 => to_slv(opcode_type, 16#DE#),
      1926 => to_slv(opcode_type, 16#04#),
      1927 => to_slv(opcode_type, 16#0B#),
      1928 => to_slv(opcode_type, 16#08#),
      1929 => to_slv(opcode_type, 16#09#),
      1930 => to_slv(opcode_type, 16#0D#),
      1931 => to_slv(opcode_type, 16#29#),
      1932 => to_slv(opcode_type, 16#08#),
      1933 => to_slv(opcode_type, 16#0B#),
      1934 => to_slv(opcode_type, 16#0A#),
      1935 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#05#),
      1953 => to_slv(opcode_type, 16#06#),
      1954 => to_slv(opcode_type, 16#08#),
      1955 => to_slv(opcode_type, 16#04#),
      1956 => to_slv(opcode_type, 16#B8#),
      1957 => to_slv(opcode_type, 16#07#),
      1958 => to_slv(opcode_type, 16#16#),
      1959 => to_slv(opcode_type, 16#A5#),
      1960 => to_slv(opcode_type, 16#08#),
      1961 => to_slv(opcode_type, 16#06#),
      1962 => to_slv(opcode_type, 16#0A#),
      1963 => to_slv(opcode_type, 16#10#),
      1964 => to_slv(opcode_type, 16#06#),
      1965 => to_slv(opcode_type, 16#11#),
      1966 => to_slv(opcode_type, 16#0B#),
      1967 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#09#),
      1985 => to_slv(opcode_type, 16#01#),
      1986 => to_slv(opcode_type, 16#04#),
      1987 => to_slv(opcode_type, 16#02#),
      1988 => to_slv(opcode_type, 16#0F#),
      1989 => to_slv(opcode_type, 16#06#),
      1990 => to_slv(opcode_type, 16#03#),
      1991 => to_slv(opcode_type, 16#05#),
      1992 => to_slv(opcode_type, 16#0C#),
      1993 => to_slv(opcode_type, 16#07#),
      1994 => to_slv(opcode_type, 16#02#),
      1995 => to_slv(opcode_type, 16#0C#),
      1996 => to_slv(opcode_type, 16#06#),
      1997 => to_slv(opcode_type, 16#0E#),
      1998 => to_slv(opcode_type, 16#11#),
      1999 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#07#),
      2017 => to_slv(opcode_type, 16#04#),
      2018 => to_slv(opcode_type, 16#09#),
      2019 => to_slv(opcode_type, 16#07#),
      2020 => to_slv(opcode_type, 16#0D#),
      2021 => to_slv(opcode_type, 16#1F#),
      2022 => to_slv(opcode_type, 16#01#),
      2023 => to_slv(opcode_type, 16#11#),
      2024 => to_slv(opcode_type, 16#01#),
      2025 => to_slv(opcode_type, 16#07#),
      2026 => to_slv(opcode_type, 16#04#),
      2027 => to_slv(opcode_type, 16#0D#),
      2028 => to_slv(opcode_type, 16#08#),
      2029 => to_slv(opcode_type, 16#0C#),
      2030 => to_slv(opcode_type, 16#10#),
      2031 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#03#),
      2049 => to_slv(opcode_type, 16#07#),
      2050 => to_slv(opcode_type, 16#07#),
      2051 => to_slv(opcode_type, 16#09#),
      2052 => to_slv(opcode_type, 16#11#),
      2053 => to_slv(opcode_type, 16#0B#),
      2054 => to_slv(opcode_type, 16#01#),
      2055 => to_slv(opcode_type, 16#0B#),
      2056 => to_slv(opcode_type, 16#09#),
      2057 => to_slv(opcode_type, 16#08#),
      2058 => to_slv(opcode_type, 16#0B#),
      2059 => to_slv(opcode_type, 16#2B#),
      2060 => to_slv(opcode_type, 16#07#),
      2061 => to_slv(opcode_type, 16#10#),
      2062 => to_slv(opcode_type, 16#0F#),
      2063 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#02#),
      2081 => to_slv(opcode_type, 16#06#),
      2082 => to_slv(opcode_type, 16#06#),
      2083 => to_slv(opcode_type, 16#06#),
      2084 => to_slv(opcode_type, 16#0B#),
      2085 => to_slv(opcode_type, 16#0E#),
      2086 => to_slv(opcode_type, 16#06#),
      2087 => to_slv(opcode_type, 16#0A#),
      2088 => to_slv(opcode_type, 16#0B#),
      2089 => to_slv(opcode_type, 16#09#),
      2090 => to_slv(opcode_type, 16#09#),
      2091 => to_slv(opcode_type, 16#0B#),
      2092 => to_slv(opcode_type, 16#0F#),
      2093 => to_slv(opcode_type, 16#05#),
      2094 => to_slv(opcode_type, 16#10#),
      2095 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#04#),
      2113 => to_slv(opcode_type, 16#06#),
      2114 => to_slv(opcode_type, 16#09#),
      2115 => to_slv(opcode_type, 16#09#),
      2116 => to_slv(opcode_type, 16#0F#),
      2117 => to_slv(opcode_type, 16#0B#),
      2118 => to_slv(opcode_type, 16#01#),
      2119 => to_slv(opcode_type, 16#10#),
      2120 => to_slv(opcode_type, 16#07#),
      2121 => to_slv(opcode_type, 16#06#),
      2122 => to_slv(opcode_type, 16#11#),
      2123 => to_slv(opcode_type, 16#10#),
      2124 => to_slv(opcode_type, 16#07#),
      2125 => to_slv(opcode_type, 16#55#),
      2126 => to_slv(opcode_type, 16#0D#),
      2127 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#08#),
      2146 => to_slv(opcode_type, 16#04#),
      2147 => to_slv(opcode_type, 16#02#),
      2148 => to_slv(opcode_type, 16#0E#),
      2149 => to_slv(opcode_type, 16#08#),
      2150 => to_slv(opcode_type, 16#04#),
      2151 => to_slv(opcode_type, 16#0C#),
      2152 => to_slv(opcode_type, 16#09#),
      2153 => to_slv(opcode_type, 16#0D#),
      2154 => to_slv(opcode_type, 16#0E#),
      2155 => to_slv(opcode_type, 16#07#),
      2156 => to_slv(opcode_type, 16#01#),
      2157 => to_slv(opcode_type, 16#0B#),
      2158 => to_slv(opcode_type, 16#0A#),
      2159 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#04#),
      2177 => to_slv(opcode_type, 16#09#),
      2178 => to_slv(opcode_type, 16#06#),
      2179 => to_slv(opcode_type, 16#06#),
      2180 => to_slv(opcode_type, 16#0B#),
      2181 => to_slv(opcode_type, 16#0A#),
      2182 => to_slv(opcode_type, 16#02#),
      2183 => to_slv(opcode_type, 16#0B#),
      2184 => to_slv(opcode_type, 16#06#),
      2185 => to_slv(opcode_type, 16#09#),
      2186 => to_slv(opcode_type, 16#0F#),
      2187 => to_slv(opcode_type, 16#0C#),
      2188 => to_slv(opcode_type, 16#07#),
      2189 => to_slv(opcode_type, 16#0B#),
      2190 => to_slv(opcode_type, 16#10#),
      2191 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#07#),
      2209 => to_slv(opcode_type, 16#08#),
      2210 => to_slv(opcode_type, 16#09#),
      2211 => to_slv(opcode_type, 16#07#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#10#),
      2214 => to_slv(opcode_type, 16#02#),
      2215 => to_slv(opcode_type, 16#0A#),
      2216 => to_slv(opcode_type, 16#08#),
      2217 => to_slv(opcode_type, 16#02#),
      2218 => to_slv(opcode_type, 16#0A#),
      2219 => to_slv(opcode_type, 16#08#),
      2220 => to_slv(opcode_type, 16#0D#),
      2221 => to_slv(opcode_type, 16#3F#),
      2222 => to_slv(opcode_type, 16#0B#),
      2223 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#01#),
      2241 => to_slv(opcode_type, 16#07#),
      2242 => to_slv(opcode_type, 16#09#),
      2243 => to_slv(opcode_type, 16#08#),
      2244 => to_slv(opcode_type, 16#0A#),
      2245 => to_slv(opcode_type, 16#0F#),
      2246 => to_slv(opcode_type, 16#05#),
      2247 => to_slv(opcode_type, 16#0C#),
      2248 => to_slv(opcode_type, 16#07#),
      2249 => to_slv(opcode_type, 16#06#),
      2250 => to_slv(opcode_type, 16#10#),
      2251 => to_slv(opcode_type, 16#0E#),
      2252 => to_slv(opcode_type, 16#06#),
      2253 => to_slv(opcode_type, 16#0C#),
      2254 => to_slv(opcode_type, 16#0F#),
      2255 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#01#),
      2273 => to_slv(opcode_type, 16#08#),
      2274 => to_slv(opcode_type, 16#07#),
      2275 => to_slv(opcode_type, 16#03#),
      2276 => to_slv(opcode_type, 16#0B#),
      2277 => to_slv(opcode_type, 16#09#),
      2278 => to_slv(opcode_type, 16#10#),
      2279 => to_slv(opcode_type, 16#0A#),
      2280 => to_slv(opcode_type, 16#07#),
      2281 => to_slv(opcode_type, 16#08#),
      2282 => to_slv(opcode_type, 16#0F#),
      2283 => to_slv(opcode_type, 16#0E#),
      2284 => to_slv(opcode_type, 16#08#),
      2285 => to_slv(opcode_type, 16#0A#),
      2286 => to_slv(opcode_type, 16#0F#),
      2287 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#01#),
      2305 => to_slv(opcode_type, 16#06#),
      2306 => to_slv(opcode_type, 16#07#),
      2307 => to_slv(opcode_type, 16#01#),
      2308 => to_slv(opcode_type, 16#10#),
      2309 => to_slv(opcode_type, 16#07#),
      2310 => to_slv(opcode_type, 16#0D#),
      2311 => to_slv(opcode_type, 16#0C#),
      2312 => to_slv(opcode_type, 16#07#),
      2313 => to_slv(opcode_type, 16#09#),
      2314 => to_slv(opcode_type, 16#0A#),
      2315 => to_slv(opcode_type, 16#0D#),
      2316 => to_slv(opcode_type, 16#07#),
      2317 => to_slv(opcode_type, 16#0D#),
      2318 => to_slv(opcode_type, 16#10#),
      2319 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#03#),
      2337 => to_slv(opcode_type, 16#07#),
      2338 => to_slv(opcode_type, 16#09#),
      2339 => to_slv(opcode_type, 16#03#),
      2340 => to_slv(opcode_type, 16#0A#),
      2341 => to_slv(opcode_type, 16#07#),
      2342 => to_slv(opcode_type, 16#0E#),
      2343 => to_slv(opcode_type, 16#0D#),
      2344 => to_slv(opcode_type, 16#09#),
      2345 => to_slv(opcode_type, 16#08#),
      2346 => to_slv(opcode_type, 16#D3#),
      2347 => to_slv(opcode_type, 16#0A#),
      2348 => to_slv(opcode_type, 16#08#),
      2349 => to_slv(opcode_type, 16#0B#),
      2350 => to_slv(opcode_type, 16#0E#),
      2351 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#01#),
      2369 => to_slv(opcode_type, 16#07#),
      2370 => to_slv(opcode_type, 16#06#),
      2371 => to_slv(opcode_type, 16#06#),
      2372 => to_slv(opcode_type, 16#10#),
      2373 => to_slv(opcode_type, 16#5C#),
      2374 => to_slv(opcode_type, 16#03#),
      2375 => to_slv(opcode_type, 16#0C#),
      2376 => to_slv(opcode_type, 16#08#),
      2377 => to_slv(opcode_type, 16#08#),
      2378 => to_slv(opcode_type, 16#11#),
      2379 => to_slv(opcode_type, 16#0B#),
      2380 => to_slv(opcode_type, 16#06#),
      2381 => to_slv(opcode_type, 16#0A#),
      2382 => to_slv(opcode_type, 16#0D#),
      2383 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#01#),
      2402 => to_slv(opcode_type, 16#01#),
      2403 => to_slv(opcode_type, 16#06#),
      2404 => to_slv(opcode_type, 16#20#),
      2405 => to_slv(opcode_type, 16#0B#),
      2406 => to_slv(opcode_type, 16#09#),
      2407 => to_slv(opcode_type, 16#03#),
      2408 => to_slv(opcode_type, 16#01#),
      2409 => to_slv(opcode_type, 16#0F#),
      2410 => to_slv(opcode_type, 16#07#),
      2411 => to_slv(opcode_type, 16#06#),
      2412 => to_slv(opcode_type, 16#0A#),
      2413 => to_slv(opcode_type, 16#2F#),
      2414 => to_slv(opcode_type, 16#0E#),
      2415 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#07#),
      2433 => to_slv(opcode_type, 16#04#),
      2434 => to_slv(opcode_type, 16#04#),
      2435 => to_slv(opcode_type, 16#05#),
      2436 => to_slv(opcode_type, 16#0A#),
      2437 => to_slv(opcode_type, 16#09#),
      2438 => to_slv(opcode_type, 16#06#),
      2439 => to_slv(opcode_type, 16#01#),
      2440 => to_slv(opcode_type, 16#6F#),
      2441 => to_slv(opcode_type, 16#02#),
      2442 => to_slv(opcode_type, 16#0D#),
      2443 => to_slv(opcode_type, 16#02#),
      2444 => to_slv(opcode_type, 16#06#),
      2445 => to_slv(opcode_type, 16#0D#),
      2446 => to_slv(opcode_type, 16#0E#),
      2447 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#07#),
      2465 => to_slv(opcode_type, 16#02#),
      2466 => to_slv(opcode_type, 16#03#),
      2467 => to_slv(opcode_type, 16#01#),
      2468 => to_slv(opcode_type, 16#0B#),
      2469 => to_slv(opcode_type, 16#08#),
      2470 => to_slv(opcode_type, 16#04#),
      2471 => to_slv(opcode_type, 16#09#),
      2472 => to_slv(opcode_type, 16#0C#),
      2473 => to_slv(opcode_type, 16#10#),
      2474 => to_slv(opcode_type, 16#08#),
      2475 => to_slv(opcode_type, 16#02#),
      2476 => to_slv(opcode_type, 16#10#),
      2477 => to_slv(opcode_type, 16#02#),
      2478 => to_slv(opcode_type, 16#0B#),
      2479 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#01#),
      2497 => to_slv(opcode_type, 16#07#),
      2498 => to_slv(opcode_type, 16#07#),
      2499 => to_slv(opcode_type, 16#07#),
      2500 => to_slv(opcode_type, 16#0F#),
      2501 => to_slv(opcode_type, 16#11#),
      2502 => to_slv(opcode_type, 16#07#),
      2503 => to_slv(opcode_type, 16#11#),
      2504 => to_slv(opcode_type, 16#11#),
      2505 => to_slv(opcode_type, 16#08#),
      2506 => to_slv(opcode_type, 16#06#),
      2507 => to_slv(opcode_type, 16#0C#),
      2508 => to_slv(opcode_type, 16#0F#),
      2509 => to_slv(opcode_type, 16#04#),
      2510 => to_slv(opcode_type, 16#35#),
      2511 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#01#),
      2529 => to_slv(opcode_type, 16#06#),
      2530 => to_slv(opcode_type, 16#08#),
      2531 => to_slv(opcode_type, 16#09#),
      2532 => to_slv(opcode_type, 16#0E#),
      2533 => to_slv(opcode_type, 16#0F#),
      2534 => to_slv(opcode_type, 16#08#),
      2535 => to_slv(opcode_type, 16#0D#),
      2536 => to_slv(opcode_type, 16#0F#),
      2537 => to_slv(opcode_type, 16#09#),
      2538 => to_slv(opcode_type, 16#08#),
      2539 => to_slv(opcode_type, 16#6B#),
      2540 => to_slv(opcode_type, 16#10#),
      2541 => to_slv(opcode_type, 16#05#),
      2542 => to_slv(opcode_type, 16#10#),
      2543 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#05#),
      2561 => to_slv(opcode_type, 16#07#),
      2562 => to_slv(opcode_type, 16#09#),
      2563 => to_slv(opcode_type, 16#05#),
      2564 => to_slv(opcode_type, 16#0D#),
      2565 => to_slv(opcode_type, 16#09#),
      2566 => to_slv(opcode_type, 16#0B#),
      2567 => to_slv(opcode_type, 16#0B#),
      2568 => to_slv(opcode_type, 16#06#),
      2569 => to_slv(opcode_type, 16#06#),
      2570 => to_slv(opcode_type, 16#10#),
      2571 => to_slv(opcode_type, 16#0F#),
      2572 => to_slv(opcode_type, 16#09#),
      2573 => to_slv(opcode_type, 16#0E#),
      2574 => to_slv(opcode_type, 16#10#),
      2575 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#07#),
      2593 => to_slv(opcode_type, 16#02#),
      2594 => to_slv(opcode_type, 16#09#),
      2595 => to_slv(opcode_type, 16#02#),
      2596 => to_slv(opcode_type, 16#0D#),
      2597 => to_slv(opcode_type, 16#05#),
      2598 => to_slv(opcode_type, 16#0C#),
      2599 => to_slv(opcode_type, 16#07#),
      2600 => to_slv(opcode_type, 16#01#),
      2601 => to_slv(opcode_type, 16#07#),
      2602 => to_slv(opcode_type, 16#10#),
      2603 => to_slv(opcode_type, 16#11#),
      2604 => to_slv(opcode_type, 16#05#),
      2605 => to_slv(opcode_type, 16#03#),
      2606 => to_slv(opcode_type, 16#0E#),
      2607 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#05#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#09#),
      2627 => to_slv(opcode_type, 16#04#),
      2628 => to_slv(opcode_type, 16#0D#),
      2629 => to_slv(opcode_type, 16#07#),
      2630 => to_slv(opcode_type, 16#10#),
      2631 => to_slv(opcode_type, 16#11#),
      2632 => to_slv(opcode_type, 16#07#),
      2633 => to_slv(opcode_type, 16#08#),
      2634 => to_slv(opcode_type, 16#0A#),
      2635 => to_slv(opcode_type, 16#11#),
      2636 => to_slv(opcode_type, 16#07#),
      2637 => to_slv(opcode_type, 16#0F#),
      2638 => to_slv(opcode_type, 16#0D#),
      2639 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#05#),
      2657 => to_slv(opcode_type, 16#07#),
      2658 => to_slv(opcode_type, 16#07#),
      2659 => to_slv(opcode_type, 16#07#),
      2660 => to_slv(opcode_type, 16#0E#),
      2661 => to_slv(opcode_type, 16#11#),
      2662 => to_slv(opcode_type, 16#01#),
      2663 => to_slv(opcode_type, 16#A8#),
      2664 => to_slv(opcode_type, 16#07#),
      2665 => to_slv(opcode_type, 16#06#),
      2666 => to_slv(opcode_type, 16#0F#),
      2667 => to_slv(opcode_type, 16#82#),
      2668 => to_slv(opcode_type, 16#07#),
      2669 => to_slv(opcode_type, 16#0E#),
      2670 => to_slv(opcode_type, 16#0F#),
      2671 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#06#),
      2689 => to_slv(opcode_type, 16#02#),
      2690 => to_slv(opcode_type, 16#03#),
      2691 => to_slv(opcode_type, 16#06#),
      2692 => to_slv(opcode_type, 16#0E#),
      2693 => to_slv(opcode_type, 16#0B#),
      2694 => to_slv(opcode_type, 16#06#),
      2695 => to_slv(opcode_type, 16#02#),
      2696 => to_slv(opcode_type, 16#06#),
      2697 => to_slv(opcode_type, 16#0D#),
      2698 => to_slv(opcode_type, 16#0D#),
      2699 => to_slv(opcode_type, 16#08#),
      2700 => to_slv(opcode_type, 16#03#),
      2701 => to_slv(opcode_type, 16#11#),
      2702 => to_slv(opcode_type, 16#0B#),
      2703 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#07#),
      2721 => to_slv(opcode_type, 16#03#),
      2722 => to_slv(opcode_type, 16#04#),
      2723 => to_slv(opcode_type, 16#08#),
      2724 => to_slv(opcode_type, 16#11#),
      2725 => to_slv(opcode_type, 16#0D#),
      2726 => to_slv(opcode_type, 16#07#),
      2727 => to_slv(opcode_type, 16#03#),
      2728 => to_slv(opcode_type, 16#07#),
      2729 => to_slv(opcode_type, 16#0F#),
      2730 => to_slv(opcode_type, 16#11#),
      2731 => to_slv(opcode_type, 16#05#),
      2732 => to_slv(opcode_type, 16#06#),
      2733 => to_slv(opcode_type, 16#0A#),
      2734 => to_slv(opcode_type, 16#0D#),
      2735 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#05#),
      2753 => to_slv(opcode_type, 16#09#),
      2754 => to_slv(opcode_type, 16#09#),
      2755 => to_slv(opcode_type, 16#09#),
      2756 => to_slv(opcode_type, 16#0F#),
      2757 => to_slv(opcode_type, 16#0A#),
      2758 => to_slv(opcode_type, 16#01#),
      2759 => to_slv(opcode_type, 16#0C#),
      2760 => to_slv(opcode_type, 16#08#),
      2761 => to_slv(opcode_type, 16#06#),
      2762 => to_slv(opcode_type, 16#11#),
      2763 => to_slv(opcode_type, 16#0F#),
      2764 => to_slv(opcode_type, 16#06#),
      2765 => to_slv(opcode_type, 16#0F#),
      2766 => to_slv(opcode_type, 16#0B#),
      2767 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#09#),
      2785 => to_slv(opcode_type, 16#03#),
      2786 => to_slv(opcode_type, 16#03#),
      2787 => to_slv(opcode_type, 16#07#),
      2788 => to_slv(opcode_type, 16#0A#),
      2789 => to_slv(opcode_type, 16#0E#),
      2790 => to_slv(opcode_type, 16#07#),
      2791 => to_slv(opcode_type, 16#03#),
      2792 => to_slv(opcode_type, 16#02#),
      2793 => to_slv(opcode_type, 16#10#),
      2794 => to_slv(opcode_type, 16#07#),
      2795 => to_slv(opcode_type, 16#05#),
      2796 => to_slv(opcode_type, 16#0A#),
      2797 => to_slv(opcode_type, 16#01#),
      2798 => to_slv(opcode_type, 16#10#),
      2799 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#06#),
      2817 => to_slv(opcode_type, 16#02#),
      2818 => to_slv(opcode_type, 16#05#),
      2819 => to_slv(opcode_type, 16#06#),
      2820 => to_slv(opcode_type, 16#10#),
      2821 => to_slv(opcode_type, 16#0C#),
      2822 => to_slv(opcode_type, 16#09#),
      2823 => to_slv(opcode_type, 16#03#),
      2824 => to_slv(opcode_type, 16#06#),
      2825 => to_slv(opcode_type, 16#0D#),
      2826 => to_slv(opcode_type, 16#0D#),
      2827 => to_slv(opcode_type, 16#09#),
      2828 => to_slv(opcode_type, 16#02#),
      2829 => to_slv(opcode_type, 16#10#),
      2830 => to_slv(opcode_type, 16#11#),
      2831 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#07#),
      2849 => to_slv(opcode_type, 16#01#),
      2850 => to_slv(opcode_type, 16#08#),
      2851 => to_slv(opcode_type, 16#05#),
      2852 => to_slv(opcode_type, 16#0E#),
      2853 => to_slv(opcode_type, 16#04#),
      2854 => to_slv(opcode_type, 16#10#),
      2855 => to_slv(opcode_type, 16#09#),
      2856 => to_slv(opcode_type, 16#02#),
      2857 => to_slv(opcode_type, 16#05#),
      2858 => to_slv(opcode_type, 16#0F#),
      2859 => to_slv(opcode_type, 16#05#),
      2860 => to_slv(opcode_type, 16#08#),
      2861 => to_slv(opcode_type, 16#11#),
      2862 => to_slv(opcode_type, 16#0A#),
      2863 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#05#),
      2881 => to_slv(opcode_type, 16#07#),
      2882 => to_slv(opcode_type, 16#06#),
      2883 => to_slv(opcode_type, 16#08#),
      2884 => to_slv(opcode_type, 16#0D#),
      2885 => to_slv(opcode_type, 16#0E#),
      2886 => to_slv(opcode_type, 16#09#),
      2887 => to_slv(opcode_type, 16#10#),
      2888 => to_slv(opcode_type, 16#0F#),
      2889 => to_slv(opcode_type, 16#07#),
      2890 => to_slv(opcode_type, 16#04#),
      2891 => to_slv(opcode_type, 16#0E#),
      2892 => to_slv(opcode_type, 16#08#),
      2893 => to_slv(opcode_type, 16#0A#),
      2894 => to_slv(opcode_type, 16#0E#),
      2895 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#01#),
      2913 => to_slv(opcode_type, 16#06#),
      2914 => to_slv(opcode_type, 16#09#),
      2915 => to_slv(opcode_type, 16#09#),
      2916 => to_slv(opcode_type, 16#0F#),
      2917 => to_slv(opcode_type, 16#0D#),
      2918 => to_slv(opcode_type, 16#09#),
      2919 => to_slv(opcode_type, 16#0D#),
      2920 => to_slv(opcode_type, 16#0D#),
      2921 => to_slv(opcode_type, 16#08#),
      2922 => to_slv(opcode_type, 16#09#),
      2923 => to_slv(opcode_type, 16#0E#),
      2924 => to_slv(opcode_type, 16#0A#),
      2925 => to_slv(opcode_type, 16#05#),
      2926 => to_slv(opcode_type, 16#0B#),
      2927 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#07#),
      2945 => to_slv(opcode_type, 16#05#),
      2946 => to_slv(opcode_type, 16#05#),
      2947 => to_slv(opcode_type, 16#03#),
      2948 => to_slv(opcode_type, 16#0B#),
      2949 => to_slv(opcode_type, 16#06#),
      2950 => to_slv(opcode_type, 16#01#),
      2951 => to_slv(opcode_type, 16#07#),
      2952 => to_slv(opcode_type, 16#10#),
      2953 => to_slv(opcode_type, 16#0F#),
      2954 => to_slv(opcode_type, 16#09#),
      2955 => to_slv(opcode_type, 16#09#),
      2956 => to_slv(opcode_type, 16#0C#),
      2957 => to_slv(opcode_type, 16#0D#),
      2958 => to_slv(opcode_type, 16#0F#),
      2959 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#02#),
      2977 => to_slv(opcode_type, 16#08#),
      2978 => to_slv(opcode_type, 16#06#),
      2979 => to_slv(opcode_type, 16#03#),
      2980 => to_slv(opcode_type, 16#0D#),
      2981 => to_slv(opcode_type, 16#07#),
      2982 => to_slv(opcode_type, 16#0B#),
      2983 => to_slv(opcode_type, 16#0C#),
      2984 => to_slv(opcode_type, 16#09#),
      2985 => to_slv(opcode_type, 16#09#),
      2986 => to_slv(opcode_type, 16#0E#),
      2987 => to_slv(opcode_type, 16#10#),
      2988 => to_slv(opcode_type, 16#06#),
      2989 => to_slv(opcode_type, 16#0E#),
      2990 => to_slv(opcode_type, 16#10#),
      2991 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#08#),
      3009 => to_slv(opcode_type, 16#06#),
      3010 => to_slv(opcode_type, 16#09#),
      3011 => to_slv(opcode_type, 16#06#),
      3012 => to_slv(opcode_type, 16#0E#),
      3013 => to_slv(opcode_type, 16#0B#),
      3014 => to_slv(opcode_type, 16#03#),
      3015 => to_slv(opcode_type, 16#0F#),
      3016 => to_slv(opcode_type, 16#01#),
      3017 => to_slv(opcode_type, 16#02#),
      3018 => to_slv(opcode_type, 16#0F#),
      3019 => to_slv(opcode_type, 16#01#),
      3020 => to_slv(opcode_type, 16#05#),
      3021 => to_slv(opcode_type, 16#05#),
      3022 => to_slv(opcode_type, 16#0A#),
      3023 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#04#),
      3041 => to_slv(opcode_type, 16#06#),
      3042 => to_slv(opcode_type, 16#09#),
      3043 => to_slv(opcode_type, 16#09#),
      3044 => to_slv(opcode_type, 16#0E#),
      3045 => to_slv(opcode_type, 16#11#),
      3046 => to_slv(opcode_type, 16#02#),
      3047 => to_slv(opcode_type, 16#0B#),
      3048 => to_slv(opcode_type, 16#08#),
      3049 => to_slv(opcode_type, 16#09#),
      3050 => to_slv(opcode_type, 16#0A#),
      3051 => to_slv(opcode_type, 16#10#),
      3052 => to_slv(opcode_type, 16#06#),
      3053 => to_slv(opcode_type, 16#11#),
      3054 => to_slv(opcode_type, 16#10#),
      3055 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#05#),
      3073 => to_slv(opcode_type, 16#06#),
      3074 => to_slv(opcode_type, 16#07#),
      3075 => to_slv(opcode_type, 16#08#),
      3076 => to_slv(opcode_type, 16#11#),
      3077 => to_slv(opcode_type, 16#25#),
      3078 => to_slv(opcode_type, 16#08#),
      3079 => to_slv(opcode_type, 16#0E#),
      3080 => to_slv(opcode_type, 16#0A#),
      3081 => to_slv(opcode_type, 16#09#),
      3082 => to_slv(opcode_type, 16#03#),
      3083 => to_slv(opcode_type, 16#0B#),
      3084 => to_slv(opcode_type, 16#07#),
      3085 => to_slv(opcode_type, 16#10#),
      3086 => to_slv(opcode_type, 16#74#),
      3087 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#05#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#07#),
      3107 => to_slv(opcode_type, 16#06#),
      3108 => to_slv(opcode_type, 16#11#),
      3109 => to_slv(opcode_type, 16#0E#),
      3110 => to_slv(opcode_type, 16#09#),
      3111 => to_slv(opcode_type, 16#0D#),
      3112 => to_slv(opcode_type, 16#AE#),
      3113 => to_slv(opcode_type, 16#08#),
      3114 => to_slv(opcode_type, 16#07#),
      3115 => to_slv(opcode_type, 16#0B#),
      3116 => to_slv(opcode_type, 16#0C#),
      3117 => to_slv(opcode_type, 16#01#),
      3118 => to_slv(opcode_type, 16#10#),
      3119 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#06#),
      3137 => to_slv(opcode_type, 16#01#),
      3138 => to_slv(opcode_type, 16#02#),
      3139 => to_slv(opcode_type, 16#07#),
      3140 => to_slv(opcode_type, 16#10#),
      3141 => to_slv(opcode_type, 16#0D#),
      3142 => to_slv(opcode_type, 16#09#),
      3143 => to_slv(opcode_type, 16#07#),
      3144 => to_slv(opcode_type, 16#03#),
      3145 => to_slv(opcode_type, 16#0D#),
      3146 => to_slv(opcode_type, 16#08#),
      3147 => to_slv(opcode_type, 16#11#),
      3148 => to_slv(opcode_type, 16#80#),
      3149 => to_slv(opcode_type, 16#04#),
      3150 => to_slv(opcode_type, 16#0D#),
      3151 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#05#),
      3169 => to_slv(opcode_type, 16#06#),
      3170 => to_slv(opcode_type, 16#09#),
      3171 => to_slv(opcode_type, 16#04#),
      3172 => to_slv(opcode_type, 16#0F#),
      3173 => to_slv(opcode_type, 16#07#),
      3174 => to_slv(opcode_type, 16#D3#),
      3175 => to_slv(opcode_type, 16#0A#),
      3176 => to_slv(opcode_type, 16#07#),
      3177 => to_slv(opcode_type, 16#07#),
      3178 => to_slv(opcode_type, 16#0F#),
      3179 => to_slv(opcode_type, 16#0A#),
      3180 => to_slv(opcode_type, 16#06#),
      3181 => to_slv(opcode_type, 16#0B#),
      3182 => to_slv(opcode_type, 16#11#),
      3183 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#07#),
      3201 => to_slv(opcode_type, 16#01#),
      3202 => to_slv(opcode_type, 16#01#),
      3203 => to_slv(opcode_type, 16#09#),
      3204 => to_slv(opcode_type, 16#11#),
      3205 => to_slv(opcode_type, 16#0C#),
      3206 => to_slv(opcode_type, 16#09#),
      3207 => to_slv(opcode_type, 16#09#),
      3208 => to_slv(opcode_type, 16#01#),
      3209 => to_slv(opcode_type, 16#0F#),
      3210 => to_slv(opcode_type, 16#07#),
      3211 => to_slv(opcode_type, 16#0D#),
      3212 => to_slv(opcode_type, 16#2F#),
      3213 => to_slv(opcode_type, 16#02#),
      3214 => to_slv(opcode_type, 16#0B#),
      3215 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#05#),
      3234 => to_slv(opcode_type, 16#09#),
      3235 => to_slv(opcode_type, 16#02#),
      3236 => to_slv(opcode_type, 16#0D#),
      3237 => to_slv(opcode_type, 16#04#),
      3238 => to_slv(opcode_type, 16#0A#),
      3239 => to_slv(opcode_type, 16#01#),
      3240 => to_slv(opcode_type, 16#09#),
      3241 => to_slv(opcode_type, 16#06#),
      3242 => to_slv(opcode_type, 16#0E#),
      3243 => to_slv(opcode_type, 16#11#),
      3244 => to_slv(opcode_type, 16#06#),
      3245 => to_slv(opcode_type, 16#11#),
      3246 => to_slv(opcode_type, 16#0C#),
      3247 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#03#),
      3265 => to_slv(opcode_type, 16#09#),
      3266 => to_slv(opcode_type, 16#08#),
      3267 => to_slv(opcode_type, 16#08#),
      3268 => to_slv(opcode_type, 16#0B#),
      3269 => to_slv(opcode_type, 16#71#),
      3270 => to_slv(opcode_type, 16#04#),
      3271 => to_slv(opcode_type, 16#24#),
      3272 => to_slv(opcode_type, 16#07#),
      3273 => to_slv(opcode_type, 16#06#),
      3274 => to_slv(opcode_type, 16#FE#),
      3275 => to_slv(opcode_type, 16#10#),
      3276 => to_slv(opcode_type, 16#09#),
      3277 => to_slv(opcode_type, 16#10#),
      3278 => to_slv(opcode_type, 16#14#),
      3279 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#03#),
      3297 => to_slv(opcode_type, 16#06#),
      3298 => to_slv(opcode_type, 16#06#),
      3299 => to_slv(opcode_type, 16#09#),
      3300 => to_slv(opcode_type, 16#0D#),
      3301 => to_slv(opcode_type, 16#0E#),
      3302 => to_slv(opcode_type, 16#09#),
      3303 => to_slv(opcode_type, 16#7B#),
      3304 => to_slv(opcode_type, 16#FA#),
      3305 => to_slv(opcode_type, 16#09#),
      3306 => to_slv(opcode_type, 16#07#),
      3307 => to_slv(opcode_type, 16#10#),
      3308 => to_slv(opcode_type, 16#11#),
      3309 => to_slv(opcode_type, 16#05#),
      3310 => to_slv(opcode_type, 16#11#),
      3311 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#06#),
      3329 => to_slv(opcode_type, 16#06#),
      3330 => to_slv(opcode_type, 16#05#),
      3331 => to_slv(opcode_type, 16#07#),
      3332 => to_slv(opcode_type, 16#0F#),
      3333 => to_slv(opcode_type, 16#8A#),
      3334 => to_slv(opcode_type, 16#03#),
      3335 => to_slv(opcode_type, 16#04#),
      3336 => to_slv(opcode_type, 16#0F#),
      3337 => to_slv(opcode_type, 16#08#),
      3338 => to_slv(opcode_type, 16#07#),
      3339 => to_slv(opcode_type, 16#01#),
      3340 => to_slv(opcode_type, 16#10#),
      3341 => to_slv(opcode_type, 16#2B#),
      3342 => to_slv(opcode_type, 16#9E#),
      3343 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#09#),
      3361 => to_slv(opcode_type, 16#06#),
      3362 => to_slv(opcode_type, 16#06#),
      3363 => to_slv(opcode_type, 16#01#),
      3364 => to_slv(opcode_type, 16#10#),
      3365 => to_slv(opcode_type, 16#08#),
      3366 => to_slv(opcode_type, 16#48#),
      3367 => to_slv(opcode_type, 16#0B#),
      3368 => to_slv(opcode_type, 16#04#),
      3369 => to_slv(opcode_type, 16#04#),
      3370 => to_slv(opcode_type, 16#0D#),
      3371 => to_slv(opcode_type, 16#04#),
      3372 => to_slv(opcode_type, 16#03#),
      3373 => to_slv(opcode_type, 16#04#),
      3374 => to_slv(opcode_type, 16#0B#),
      3375 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#06#),
      3393 => to_slv(opcode_type, 16#07#),
      3394 => to_slv(opcode_type, 16#08#),
      3395 => to_slv(opcode_type, 16#08#),
      3396 => to_slv(opcode_type, 16#0F#),
      3397 => to_slv(opcode_type, 16#0B#),
      3398 => to_slv(opcode_type, 16#04#),
      3399 => to_slv(opcode_type, 16#0B#),
      3400 => to_slv(opcode_type, 16#06#),
      3401 => to_slv(opcode_type, 16#08#),
      3402 => to_slv(opcode_type, 16#0F#),
      3403 => to_slv(opcode_type, 16#0A#),
      3404 => to_slv(opcode_type, 16#05#),
      3405 => to_slv(opcode_type, 16#F9#),
      3406 => to_slv(opcode_type, 16#11#),
      3407 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#02#),
      3425 => to_slv(opcode_type, 16#06#),
      3426 => to_slv(opcode_type, 16#09#),
      3427 => to_slv(opcode_type, 16#09#),
      3428 => to_slv(opcode_type, 16#0A#),
      3429 => to_slv(opcode_type, 16#0C#),
      3430 => to_slv(opcode_type, 16#01#),
      3431 => to_slv(opcode_type, 16#0E#),
      3432 => to_slv(opcode_type, 16#08#),
      3433 => to_slv(opcode_type, 16#08#),
      3434 => to_slv(opcode_type, 16#0F#),
      3435 => to_slv(opcode_type, 16#0D#),
      3436 => to_slv(opcode_type, 16#07#),
      3437 => to_slv(opcode_type, 16#0D#),
      3438 => to_slv(opcode_type, 16#10#),
      3439 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#09#),
      3457 => to_slv(opcode_type, 16#07#),
      3458 => to_slv(opcode_type, 16#08#),
      3459 => to_slv(opcode_type, 16#08#),
      3460 => to_slv(opcode_type, 16#0E#),
      3461 => to_slv(opcode_type, 16#10#),
      3462 => to_slv(opcode_type, 16#06#),
      3463 => to_slv(opcode_type, 16#0F#),
      3464 => to_slv(opcode_type, 16#0F#),
      3465 => to_slv(opcode_type, 16#03#),
      3466 => to_slv(opcode_type, 16#05#),
      3467 => to_slv(opcode_type, 16#0A#),
      3468 => to_slv(opcode_type, 16#01#),
      3469 => to_slv(opcode_type, 16#02#),
      3470 => to_slv(opcode_type, 16#0D#),
      3471 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#01#),
      3489 => to_slv(opcode_type, 16#08#),
      3490 => to_slv(opcode_type, 16#09#),
      3491 => to_slv(opcode_type, 16#01#),
      3492 => to_slv(opcode_type, 16#0D#),
      3493 => to_slv(opcode_type, 16#07#),
      3494 => to_slv(opcode_type, 16#0D#),
      3495 => to_slv(opcode_type, 16#0C#),
      3496 => to_slv(opcode_type, 16#09#),
      3497 => to_slv(opcode_type, 16#08#),
      3498 => to_slv(opcode_type, 16#0B#),
      3499 => to_slv(opcode_type, 16#0E#),
      3500 => to_slv(opcode_type, 16#07#),
      3501 => to_slv(opcode_type, 16#7C#),
      3502 => to_slv(opcode_type, 16#0B#),
      3503 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#05#),
      3521 => to_slv(opcode_type, 16#06#),
      3522 => to_slv(opcode_type, 16#08#),
      3523 => to_slv(opcode_type, 16#03#),
      3524 => to_slv(opcode_type, 16#0B#),
      3525 => to_slv(opcode_type, 16#08#),
      3526 => to_slv(opcode_type, 16#0D#),
      3527 => to_slv(opcode_type, 16#10#),
      3528 => to_slv(opcode_type, 16#08#),
      3529 => to_slv(opcode_type, 16#09#),
      3530 => to_slv(opcode_type, 16#0D#),
      3531 => to_slv(opcode_type, 16#0E#),
      3532 => to_slv(opcode_type, 16#06#),
      3533 => to_slv(opcode_type, 16#0B#),
      3534 => to_slv(opcode_type, 16#0E#),
      3535 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#09#),
      3553 => to_slv(opcode_type, 16#08#),
      3554 => to_slv(opcode_type, 16#03#),
      3555 => to_slv(opcode_type, 16#03#),
      3556 => to_slv(opcode_type, 16#10#),
      3557 => to_slv(opcode_type, 16#05#),
      3558 => to_slv(opcode_type, 16#03#),
      3559 => to_slv(opcode_type, 16#0D#),
      3560 => to_slv(opcode_type, 16#04#),
      3561 => to_slv(opcode_type, 16#07#),
      3562 => to_slv(opcode_type, 16#09#),
      3563 => to_slv(opcode_type, 16#10#),
      3564 => to_slv(opcode_type, 16#11#),
      3565 => to_slv(opcode_type, 16#05#),
      3566 => to_slv(opcode_type, 16#0F#),
      3567 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#02#),
      3585 => to_slv(opcode_type, 16#07#),
      3586 => to_slv(opcode_type, 16#07#),
      3587 => to_slv(opcode_type, 16#05#),
      3588 => to_slv(opcode_type, 16#0D#),
      3589 => to_slv(opcode_type, 16#09#),
      3590 => to_slv(opcode_type, 16#0A#),
      3591 => to_slv(opcode_type, 16#D9#),
      3592 => to_slv(opcode_type, 16#07#),
      3593 => to_slv(opcode_type, 16#06#),
      3594 => to_slv(opcode_type, 16#0D#),
      3595 => to_slv(opcode_type, 16#0A#),
      3596 => to_slv(opcode_type, 16#09#),
      3597 => to_slv(opcode_type, 16#0B#),
      3598 => to_slv(opcode_type, 16#11#),
      3599 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#02#),
      3617 => to_slv(opcode_type, 16#08#),
      3618 => to_slv(opcode_type, 16#07#),
      3619 => to_slv(opcode_type, 16#05#),
      3620 => to_slv(opcode_type, 16#0B#),
      3621 => to_slv(opcode_type, 16#07#),
      3622 => to_slv(opcode_type, 16#0C#),
      3623 => to_slv(opcode_type, 16#11#),
      3624 => to_slv(opcode_type, 16#06#),
      3625 => to_slv(opcode_type, 16#08#),
      3626 => to_slv(opcode_type, 16#11#),
      3627 => to_slv(opcode_type, 16#44#),
      3628 => to_slv(opcode_type, 16#09#),
      3629 => to_slv(opcode_type, 16#10#),
      3630 => to_slv(opcode_type, 16#11#),
      3631 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#09#),
      3649 => to_slv(opcode_type, 16#07#),
      3650 => to_slv(opcode_type, 16#02#),
      3651 => to_slv(opcode_type, 16#07#),
      3652 => to_slv(opcode_type, 16#10#),
      3653 => to_slv(opcode_type, 16#0D#),
      3654 => to_slv(opcode_type, 16#03#),
      3655 => to_slv(opcode_type, 16#06#),
      3656 => to_slv(opcode_type, 16#0E#),
      3657 => to_slv(opcode_type, 16#0A#),
      3658 => to_slv(opcode_type, 16#07#),
      3659 => to_slv(opcode_type, 16#08#),
      3660 => to_slv(opcode_type, 16#0B#),
      3661 => to_slv(opcode_type, 16#95#),
      3662 => to_slv(opcode_type, 16#11#),
      3663 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#02#),
      3681 => to_slv(opcode_type, 16#08#),
      3682 => to_slv(opcode_type, 16#07#),
      3683 => to_slv(opcode_type, 16#03#),
      3684 => to_slv(opcode_type, 16#0A#),
      3685 => to_slv(opcode_type, 16#06#),
      3686 => to_slv(opcode_type, 16#0A#),
      3687 => to_slv(opcode_type, 16#0F#),
      3688 => to_slv(opcode_type, 16#07#),
      3689 => to_slv(opcode_type, 16#07#),
      3690 => to_slv(opcode_type, 16#11#),
      3691 => to_slv(opcode_type, 16#11#),
      3692 => to_slv(opcode_type, 16#06#),
      3693 => to_slv(opcode_type, 16#E0#),
      3694 => to_slv(opcode_type, 16#10#),
      3695 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#06#),
      3713 => to_slv(opcode_type, 16#08#),
      3714 => to_slv(opcode_type, 16#08#),
      3715 => to_slv(opcode_type, 16#01#),
      3716 => to_slv(opcode_type, 16#9C#),
      3717 => to_slv(opcode_type, 16#02#),
      3718 => to_slv(opcode_type, 16#0A#),
      3719 => to_slv(opcode_type, 16#03#),
      3720 => to_slv(opcode_type, 16#08#),
      3721 => to_slv(opcode_type, 16#0D#),
      3722 => to_slv(opcode_type, 16#0B#),
      3723 => to_slv(opcode_type, 16#08#),
      3724 => to_slv(opcode_type, 16#04#),
      3725 => to_slv(opcode_type, 16#0E#),
      3726 => to_slv(opcode_type, 16#10#),
      3727 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#05#),
      3745 => to_slv(opcode_type, 16#06#),
      3746 => to_slv(opcode_type, 16#06#),
      3747 => to_slv(opcode_type, 16#07#),
      3748 => to_slv(opcode_type, 16#0B#),
      3749 => to_slv(opcode_type, 16#0D#),
      3750 => to_slv(opcode_type, 16#01#),
      3751 => to_slv(opcode_type, 16#0B#),
      3752 => to_slv(opcode_type, 16#07#),
      3753 => to_slv(opcode_type, 16#08#),
      3754 => to_slv(opcode_type, 16#10#),
      3755 => to_slv(opcode_type, 16#F0#),
      3756 => to_slv(opcode_type, 16#07#),
      3757 => to_slv(opcode_type, 16#0E#),
      3758 => to_slv(opcode_type, 16#0C#),
      3759 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#05#),
      3777 => to_slv(opcode_type, 16#09#),
      3778 => to_slv(opcode_type, 16#06#),
      3779 => to_slv(opcode_type, 16#03#),
      3780 => to_slv(opcode_type, 16#0F#),
      3781 => to_slv(opcode_type, 16#09#),
      3782 => to_slv(opcode_type, 16#0B#),
      3783 => to_slv(opcode_type, 16#0D#),
      3784 => to_slv(opcode_type, 16#06#),
      3785 => to_slv(opcode_type, 16#09#),
      3786 => to_slv(opcode_type, 16#0C#),
      3787 => to_slv(opcode_type, 16#0D#),
      3788 => to_slv(opcode_type, 16#07#),
      3789 => to_slv(opcode_type, 16#0B#),
      3790 => to_slv(opcode_type, 16#10#),
      3791 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#05#),
      3809 => to_slv(opcode_type, 16#08#),
      3810 => to_slv(opcode_type, 16#06#),
      3811 => to_slv(opcode_type, 16#05#),
      3812 => to_slv(opcode_type, 16#0C#),
      3813 => to_slv(opcode_type, 16#09#),
      3814 => to_slv(opcode_type, 16#0E#),
      3815 => to_slv(opcode_type, 16#0B#),
      3816 => to_slv(opcode_type, 16#06#),
      3817 => to_slv(opcode_type, 16#08#),
      3818 => to_slv(opcode_type, 16#0A#),
      3819 => to_slv(opcode_type, 16#0E#),
      3820 => to_slv(opcode_type, 16#06#),
      3821 => to_slv(opcode_type, 16#0A#),
      3822 => to_slv(opcode_type, 16#10#),
      3823 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#02#),
      3841 => to_slv(opcode_type, 16#09#),
      3842 => to_slv(opcode_type, 16#06#),
      3843 => to_slv(opcode_type, 16#03#),
      3844 => to_slv(opcode_type, 16#10#),
      3845 => to_slv(opcode_type, 16#06#),
      3846 => to_slv(opcode_type, 16#0A#),
      3847 => to_slv(opcode_type, 16#0D#),
      3848 => to_slv(opcode_type, 16#06#),
      3849 => to_slv(opcode_type, 16#06#),
      3850 => to_slv(opcode_type, 16#0C#),
      3851 => to_slv(opcode_type, 16#0F#),
      3852 => to_slv(opcode_type, 16#06#),
      3853 => to_slv(opcode_type, 16#0C#),
      3854 => to_slv(opcode_type, 16#0E#),
      3855 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#01#),
      3873 => to_slv(opcode_type, 16#09#),
      3874 => to_slv(opcode_type, 16#07#),
      3875 => to_slv(opcode_type, 16#04#),
      3876 => to_slv(opcode_type, 16#0F#),
      3877 => to_slv(opcode_type, 16#07#),
      3878 => to_slv(opcode_type, 16#0A#),
      3879 => to_slv(opcode_type, 16#0A#),
      3880 => to_slv(opcode_type, 16#08#),
      3881 => to_slv(opcode_type, 16#07#),
      3882 => to_slv(opcode_type, 16#11#),
      3883 => to_slv(opcode_type, 16#11#),
      3884 => to_slv(opcode_type, 16#07#),
      3885 => to_slv(opcode_type, 16#0E#),
      3886 => to_slv(opcode_type, 16#10#),
      3887 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#02#),
      3905 => to_slv(opcode_type, 16#07#),
      3906 => to_slv(opcode_type, 16#06#),
      3907 => to_slv(opcode_type, 16#04#),
      3908 => to_slv(opcode_type, 16#0E#),
      3909 => to_slv(opcode_type, 16#07#),
      3910 => to_slv(opcode_type, 16#11#),
      3911 => to_slv(opcode_type, 16#11#),
      3912 => to_slv(opcode_type, 16#06#),
      3913 => to_slv(opcode_type, 16#07#),
      3914 => to_slv(opcode_type, 16#11#),
      3915 => to_slv(opcode_type, 16#B1#),
      3916 => to_slv(opcode_type, 16#06#),
      3917 => to_slv(opcode_type, 16#0D#),
      3918 => to_slv(opcode_type, 16#0E#),
      3919 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#07#),
      3937 => to_slv(opcode_type, 16#04#),
      3938 => to_slv(opcode_type, 16#09#),
      3939 => to_slv(opcode_type, 16#09#),
      3940 => to_slv(opcode_type, 16#11#),
      3941 => to_slv(opcode_type, 16#0F#),
      3942 => to_slv(opcode_type, 16#09#),
      3943 => to_slv(opcode_type, 16#10#),
      3944 => to_slv(opcode_type, 16#10#),
      3945 => to_slv(opcode_type, 16#08#),
      3946 => to_slv(opcode_type, 16#01#),
      3947 => to_slv(opcode_type, 16#06#),
      3948 => to_slv(opcode_type, 16#10#),
      3949 => to_slv(opcode_type, 16#0E#),
      3950 => to_slv(opcode_type, 16#0E#),
      3951 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#09#),
      3969 => to_slv(opcode_type, 16#07#),
      3970 => to_slv(opcode_type, 16#06#),
      3971 => to_slv(opcode_type, 16#08#),
      3972 => to_slv(opcode_type, 16#0A#),
      3973 => to_slv(opcode_type, 16#0D#),
      3974 => to_slv(opcode_type, 16#03#),
      3975 => to_slv(opcode_type, 16#8D#),
      3976 => to_slv(opcode_type, 16#08#),
      3977 => to_slv(opcode_type, 16#09#),
      3978 => to_slv(opcode_type, 16#0F#),
      3979 => to_slv(opcode_type, 16#4F#),
      3980 => to_slv(opcode_type, 16#02#),
      3981 => to_slv(opcode_type, 16#0F#),
      3982 => to_slv(opcode_type, 16#10#),
      3983 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#06#),
      4001 => to_slv(opcode_type, 16#08#),
      4002 => to_slv(opcode_type, 16#02#),
      4003 => to_slv(opcode_type, 16#06#),
      4004 => to_slv(opcode_type, 16#11#),
      4005 => to_slv(opcode_type, 16#0A#),
      4006 => to_slv(opcode_type, 16#03#),
      4007 => to_slv(opcode_type, 16#09#),
      4008 => to_slv(opcode_type, 16#0F#),
      4009 => to_slv(opcode_type, 16#0D#),
      4010 => to_slv(opcode_type, 16#01#),
      4011 => to_slv(opcode_type, 16#01#),
      4012 => to_slv(opcode_type, 16#09#),
      4013 => to_slv(opcode_type, 16#0F#),
      4014 => to_slv(opcode_type, 16#0C#),
      4015 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#06#),
      4033 => to_slv(opcode_type, 16#01#),
      4034 => to_slv(opcode_type, 16#05#),
      4035 => to_slv(opcode_type, 16#09#),
      4036 => to_slv(opcode_type, 16#0D#),
      4037 => to_slv(opcode_type, 16#0C#),
      4038 => to_slv(opcode_type, 16#09#),
      4039 => to_slv(opcode_type, 16#02#),
      4040 => to_slv(opcode_type, 16#01#),
      4041 => to_slv(opcode_type, 16#0A#),
      4042 => to_slv(opcode_type, 16#09#),
      4043 => to_slv(opcode_type, 16#01#),
      4044 => to_slv(opcode_type, 16#0B#),
      4045 => to_slv(opcode_type, 16#02#),
      4046 => to_slv(opcode_type, 16#0F#),
      4047 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#05#),
      4065 => to_slv(opcode_type, 16#07#),
      4066 => to_slv(opcode_type, 16#06#),
      4067 => to_slv(opcode_type, 16#09#),
      4068 => to_slv(opcode_type, 16#0E#),
      4069 => to_slv(opcode_type, 16#11#),
      4070 => to_slv(opcode_type, 16#04#),
      4071 => to_slv(opcode_type, 16#0E#),
      4072 => to_slv(opcode_type, 16#06#),
      4073 => to_slv(opcode_type, 16#07#),
      4074 => to_slv(opcode_type, 16#0C#),
      4075 => to_slv(opcode_type, 16#A2#),
      4076 => to_slv(opcode_type, 16#09#),
      4077 => to_slv(opcode_type, 16#0C#),
      4078 => to_slv(opcode_type, 16#0B#),
      4079 to 4095 => (others => '0')
  ),

    -- Bin `16`...
    15 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#03#),
      1 => to_slv(opcode_type, 16#07#),
      2 => to_slv(opcode_type, 16#08#),
      3 => to_slv(opcode_type, 16#06#),
      4 => to_slv(opcode_type, 16#F9#),
      5 => to_slv(opcode_type, 16#0C#),
      6 => to_slv(opcode_type, 16#06#),
      7 => to_slv(opcode_type, 16#A1#),
      8 => to_slv(opcode_type, 16#11#),
      9 => to_slv(opcode_type, 16#09#),
      10 => to_slv(opcode_type, 16#07#),
      11 => to_slv(opcode_type, 16#0B#),
      12 => to_slv(opcode_type, 16#0E#),
      13 => to_slv(opcode_type, 16#09#),
      14 => to_slv(opcode_type, 16#0E#),
      15 => to_slv(opcode_type, 16#0E#),
      16 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#08#),
      33 => to_slv(opcode_type, 16#02#),
      34 => to_slv(opcode_type, 16#09#),
      35 => to_slv(opcode_type, 16#06#),
      36 => to_slv(opcode_type, 16#0B#),
      37 => to_slv(opcode_type, 16#0D#),
      38 => to_slv(opcode_type, 16#07#),
      39 => to_slv(opcode_type, 16#0F#),
      40 => to_slv(opcode_type, 16#7F#),
      41 => to_slv(opcode_type, 16#02#),
      42 => to_slv(opcode_type, 16#09#),
      43 => to_slv(opcode_type, 16#07#),
      44 => to_slv(opcode_type, 16#72#),
      45 => to_slv(opcode_type, 16#0B#),
      46 => to_slv(opcode_type, 16#05#),
      47 => to_slv(opcode_type, 16#11#),
      48 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#06#),
      65 => to_slv(opcode_type, 16#07#),
      66 => to_slv(opcode_type, 16#06#),
      67 => to_slv(opcode_type, 16#01#),
      68 => to_slv(opcode_type, 16#0A#),
      69 => to_slv(opcode_type, 16#05#),
      70 => to_slv(opcode_type, 16#11#),
      71 => to_slv(opcode_type, 16#01#),
      72 => to_slv(opcode_type, 16#07#),
      73 => to_slv(opcode_type, 16#0E#),
      74 => to_slv(opcode_type, 16#0C#),
      75 => to_slv(opcode_type, 16#08#),
      76 => to_slv(opcode_type, 16#07#),
      77 => to_slv(opcode_type, 16#F4#),
      78 => to_slv(opcode_type, 16#0E#),
      79 => to_slv(opcode_type, 16#0B#),
      80 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#07#),
      97 => to_slv(opcode_type, 16#03#),
      98 => to_slv(opcode_type, 16#03#),
      99 => to_slv(opcode_type, 16#03#),
      100 => to_slv(opcode_type, 16#0C#),
      101 => to_slv(opcode_type, 16#07#),
      102 => to_slv(opcode_type, 16#06#),
      103 => to_slv(opcode_type, 16#04#),
      104 => to_slv(opcode_type, 16#0A#),
      105 => to_slv(opcode_type, 16#04#),
      106 => to_slv(opcode_type, 16#0F#),
      107 => to_slv(opcode_type, 16#09#),
      108 => to_slv(opcode_type, 16#06#),
      109 => to_slv(opcode_type, 16#10#),
      110 => to_slv(opcode_type, 16#0E#),
      111 => to_slv(opcode_type, 16#0C#),
      112 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#07#),
      129 => to_slv(opcode_type, 16#05#),
      130 => to_slv(opcode_type, 16#02#),
      131 => to_slv(opcode_type, 16#09#),
      132 => to_slv(opcode_type, 16#11#),
      133 => to_slv(opcode_type, 16#0A#),
      134 => to_slv(opcode_type, 16#09#),
      135 => to_slv(opcode_type, 16#03#),
      136 => to_slv(opcode_type, 16#06#),
      137 => to_slv(opcode_type, 16#0D#),
      138 => to_slv(opcode_type, 16#11#),
      139 => to_slv(opcode_type, 16#07#),
      140 => to_slv(opcode_type, 16#09#),
      141 => to_slv(opcode_type, 16#0A#),
      142 => to_slv(opcode_type, 16#0D#),
      143 => to_slv(opcode_type, 16#0B#),
      144 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#04#),
      161 => to_slv(opcode_type, 16#06#),
      162 => to_slv(opcode_type, 16#07#),
      163 => to_slv(opcode_type, 16#08#),
      164 => to_slv(opcode_type, 16#0C#),
      165 => to_slv(opcode_type, 16#11#),
      166 => to_slv(opcode_type, 16#07#),
      167 => to_slv(opcode_type, 16#0E#),
      168 => to_slv(opcode_type, 16#0A#),
      169 => to_slv(opcode_type, 16#06#),
      170 => to_slv(opcode_type, 16#06#),
      171 => to_slv(opcode_type, 16#0B#),
      172 => to_slv(opcode_type, 16#0B#),
      173 => to_slv(opcode_type, 16#06#),
      174 => to_slv(opcode_type, 16#BD#),
      175 => to_slv(opcode_type, 16#0A#),
      176 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#01#),
      193 => to_slv(opcode_type, 16#07#),
      194 => to_slv(opcode_type, 16#06#),
      195 => to_slv(opcode_type, 16#09#),
      196 => to_slv(opcode_type, 16#0F#),
      197 => to_slv(opcode_type, 16#0F#),
      198 => to_slv(opcode_type, 16#09#),
      199 => to_slv(opcode_type, 16#0A#),
      200 => to_slv(opcode_type, 16#0B#),
      201 => to_slv(opcode_type, 16#07#),
      202 => to_slv(opcode_type, 16#09#),
      203 => to_slv(opcode_type, 16#0B#),
      204 => to_slv(opcode_type, 16#0D#),
      205 => to_slv(opcode_type, 16#09#),
      206 => to_slv(opcode_type, 16#0D#),
      207 => to_slv(opcode_type, 16#10#),
      208 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#02#),
      225 => to_slv(opcode_type, 16#07#),
      226 => to_slv(opcode_type, 16#06#),
      227 => to_slv(opcode_type, 16#07#),
      228 => to_slv(opcode_type, 16#0F#),
      229 => to_slv(opcode_type, 16#0D#),
      230 => to_slv(opcode_type, 16#09#),
      231 => to_slv(opcode_type, 16#10#),
      232 => to_slv(opcode_type, 16#3D#),
      233 => to_slv(opcode_type, 16#08#),
      234 => to_slv(opcode_type, 16#07#),
      235 => to_slv(opcode_type, 16#0C#),
      236 => to_slv(opcode_type, 16#C7#),
      237 => to_slv(opcode_type, 16#08#),
      238 => to_slv(opcode_type, 16#11#),
      239 => to_slv(opcode_type, 16#0F#),
      240 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#04#),
      257 => to_slv(opcode_type, 16#09#),
      258 => to_slv(opcode_type, 16#08#),
      259 => to_slv(opcode_type, 16#08#),
      260 => to_slv(opcode_type, 16#0B#),
      261 => to_slv(opcode_type, 16#0F#),
      262 => to_slv(opcode_type, 16#09#),
      263 => to_slv(opcode_type, 16#10#),
      264 => to_slv(opcode_type, 16#0C#),
      265 => to_slv(opcode_type, 16#07#),
      266 => to_slv(opcode_type, 16#06#),
      267 => to_slv(opcode_type, 16#0C#),
      268 => to_slv(opcode_type, 16#0B#),
      269 => to_slv(opcode_type, 16#07#),
      270 => to_slv(opcode_type, 16#0E#),
      271 => to_slv(opcode_type, 16#0C#),
      272 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#01#),
      289 => to_slv(opcode_type, 16#07#),
      290 => to_slv(opcode_type, 16#09#),
      291 => to_slv(opcode_type, 16#09#),
      292 => to_slv(opcode_type, 16#0F#),
      293 => to_slv(opcode_type, 16#BC#),
      294 => to_slv(opcode_type, 16#09#),
      295 => to_slv(opcode_type, 16#0A#),
      296 => to_slv(opcode_type, 16#0B#),
      297 => to_slv(opcode_type, 16#06#),
      298 => to_slv(opcode_type, 16#06#),
      299 => to_slv(opcode_type, 16#0B#),
      300 => to_slv(opcode_type, 16#0E#),
      301 => to_slv(opcode_type, 16#08#),
      302 => to_slv(opcode_type, 16#0B#),
      303 => to_slv(opcode_type, 16#90#),
      304 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#05#),
      321 => to_slv(opcode_type, 16#07#),
      322 => to_slv(opcode_type, 16#06#),
      323 => to_slv(opcode_type, 16#08#),
      324 => to_slv(opcode_type, 16#0A#),
      325 => to_slv(opcode_type, 16#10#),
      326 => to_slv(opcode_type, 16#08#),
      327 => to_slv(opcode_type, 16#0E#),
      328 => to_slv(opcode_type, 16#0D#),
      329 => to_slv(opcode_type, 16#07#),
      330 => to_slv(opcode_type, 16#06#),
      331 => to_slv(opcode_type, 16#0A#),
      332 => to_slv(opcode_type, 16#0F#),
      333 => to_slv(opcode_type, 16#09#),
      334 => to_slv(opcode_type, 16#0F#),
      335 => to_slv(opcode_type, 16#11#),
      336 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#08#),
      353 => to_slv(opcode_type, 16#09#),
      354 => to_slv(opcode_type, 16#01#),
      355 => to_slv(opcode_type, 16#02#),
      356 => to_slv(opcode_type, 16#10#),
      357 => to_slv(opcode_type, 16#09#),
      358 => to_slv(opcode_type, 16#08#),
      359 => to_slv(opcode_type, 16#0B#),
      360 => to_slv(opcode_type, 16#10#),
      361 => to_slv(opcode_type, 16#05#),
      362 => to_slv(opcode_type, 16#11#),
      363 => to_slv(opcode_type, 16#08#),
      364 => to_slv(opcode_type, 16#02#),
      365 => to_slv(opcode_type, 16#05#),
      366 => to_slv(opcode_type, 16#0B#),
      367 => to_slv(opcode_type, 16#10#),
      368 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#07#),
      385 => to_slv(opcode_type, 16#01#),
      386 => to_slv(opcode_type, 16#08#),
      387 => to_slv(opcode_type, 16#02#),
      388 => to_slv(opcode_type, 16#0F#),
      389 => to_slv(opcode_type, 16#06#),
      390 => to_slv(opcode_type, 16#11#),
      391 => to_slv(opcode_type, 16#10#),
      392 => to_slv(opcode_type, 16#01#),
      393 => to_slv(opcode_type, 16#08#),
      394 => to_slv(opcode_type, 16#09#),
      395 => to_slv(opcode_type, 16#0C#),
      396 => to_slv(opcode_type, 16#A4#),
      397 => to_slv(opcode_type, 16#09#),
      398 => to_slv(opcode_type, 16#10#),
      399 => to_slv(opcode_type, 16#0C#),
      400 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#09#),
      417 => to_slv(opcode_type, 16#07#),
      418 => to_slv(opcode_type, 16#08#),
      419 => to_slv(opcode_type, 16#01#),
      420 => to_slv(opcode_type, 16#0D#),
      421 => to_slv(opcode_type, 16#06#),
      422 => to_slv(opcode_type, 16#0A#),
      423 => to_slv(opcode_type, 16#0F#),
      424 => to_slv(opcode_type, 16#01#),
      425 => to_slv(opcode_type, 16#01#),
      426 => to_slv(opcode_type, 16#0F#),
      427 => to_slv(opcode_type, 16#02#),
      428 => to_slv(opcode_type, 16#06#),
      429 => to_slv(opcode_type, 16#01#),
      430 => to_slv(opcode_type, 16#10#),
      431 => to_slv(opcode_type, 16#0A#),
      432 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#02#),
      449 => to_slv(opcode_type, 16#09#),
      450 => to_slv(opcode_type, 16#09#),
      451 => to_slv(opcode_type, 16#06#),
      452 => to_slv(opcode_type, 16#0E#),
      453 => to_slv(opcode_type, 16#10#),
      454 => to_slv(opcode_type, 16#06#),
      455 => to_slv(opcode_type, 16#10#),
      456 => to_slv(opcode_type, 16#0F#),
      457 => to_slv(opcode_type, 16#06#),
      458 => to_slv(opcode_type, 16#08#),
      459 => to_slv(opcode_type, 16#94#),
      460 => to_slv(opcode_type, 16#0F#),
      461 => to_slv(opcode_type, 16#09#),
      462 => to_slv(opcode_type, 16#0A#),
      463 => to_slv(opcode_type, 16#A6#),
      464 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#04#),
      481 => to_slv(opcode_type, 16#08#),
      482 => to_slv(opcode_type, 16#07#),
      483 => to_slv(opcode_type, 16#08#),
      484 => to_slv(opcode_type, 16#0E#),
      485 => to_slv(opcode_type, 16#0B#),
      486 => to_slv(opcode_type, 16#07#),
      487 => to_slv(opcode_type, 16#0A#),
      488 => to_slv(opcode_type, 16#0C#),
      489 => to_slv(opcode_type, 16#07#),
      490 => to_slv(opcode_type, 16#08#),
      491 => to_slv(opcode_type, 16#24#),
      492 => to_slv(opcode_type, 16#10#),
      493 => to_slv(opcode_type, 16#07#),
      494 => to_slv(opcode_type, 16#B4#),
      495 => to_slv(opcode_type, 16#11#),
      496 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#08#),
      513 => to_slv(opcode_type, 16#07#),
      514 => to_slv(opcode_type, 16#08#),
      515 => to_slv(opcode_type, 16#09#),
      516 => to_slv(opcode_type, 16#0B#),
      517 => to_slv(opcode_type, 16#11#),
      518 => to_slv(opcode_type, 16#06#),
      519 => to_slv(opcode_type, 16#11#),
      520 => to_slv(opcode_type, 16#0B#),
      521 => to_slv(opcode_type, 16#04#),
      522 => to_slv(opcode_type, 16#02#),
      523 => to_slv(opcode_type, 16#0C#),
      524 => to_slv(opcode_type, 16#08#),
      525 => to_slv(opcode_type, 16#01#),
      526 => to_slv(opcode_type, 16#11#),
      527 => to_slv(opcode_type, 16#0C#),
      528 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#06#),
      545 => to_slv(opcode_type, 16#08#),
      546 => to_slv(opcode_type, 16#05#),
      547 => to_slv(opcode_type, 16#02#),
      548 => to_slv(opcode_type, 16#36#),
      549 => to_slv(opcode_type, 16#09#),
      550 => to_slv(opcode_type, 16#06#),
      551 => to_slv(opcode_type, 16#0D#),
      552 => to_slv(opcode_type, 16#0F#),
      553 => to_slv(opcode_type, 16#07#),
      554 => to_slv(opcode_type, 16#0E#),
      555 => to_slv(opcode_type, 16#0E#),
      556 => to_slv(opcode_type, 16#04#),
      557 => to_slv(opcode_type, 16#08#),
      558 => to_slv(opcode_type, 16#0B#),
      559 => to_slv(opcode_type, 16#10#),
      560 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#07#),
      577 => to_slv(opcode_type, 16#09#),
      578 => to_slv(opcode_type, 16#07#),
      579 => to_slv(opcode_type, 16#08#),
      580 => to_slv(opcode_type, 16#C1#),
      581 => to_slv(opcode_type, 16#11#),
      582 => to_slv(opcode_type, 16#08#),
      583 => to_slv(opcode_type, 16#0C#),
      584 => to_slv(opcode_type, 16#0F#),
      585 => to_slv(opcode_type, 16#01#),
      586 => to_slv(opcode_type, 16#08#),
      587 => to_slv(opcode_type, 16#0F#),
      588 => to_slv(opcode_type, 16#0B#),
      589 => to_slv(opcode_type, 16#08#),
      590 => to_slv(opcode_type, 16#0E#),
      591 => to_slv(opcode_type, 16#B9#),
      592 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#05#),
      609 => to_slv(opcode_type, 16#09#),
      610 => to_slv(opcode_type, 16#07#),
      611 => to_slv(opcode_type, 16#08#),
      612 => to_slv(opcode_type, 16#BB#),
      613 => to_slv(opcode_type, 16#0A#),
      614 => to_slv(opcode_type, 16#09#),
      615 => to_slv(opcode_type, 16#0F#),
      616 => to_slv(opcode_type, 16#10#),
      617 => to_slv(opcode_type, 16#08#),
      618 => to_slv(opcode_type, 16#09#),
      619 => to_slv(opcode_type, 16#0A#),
      620 => to_slv(opcode_type, 16#0E#),
      621 => to_slv(opcode_type, 16#08#),
      622 => to_slv(opcode_type, 16#10#),
      623 => to_slv(opcode_type, 16#0B#),
      624 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#03#),
      641 => to_slv(opcode_type, 16#06#),
      642 => to_slv(opcode_type, 16#09#),
      643 => to_slv(opcode_type, 16#07#),
      644 => to_slv(opcode_type, 16#0D#),
      645 => to_slv(opcode_type, 16#0E#),
      646 => to_slv(opcode_type, 16#09#),
      647 => to_slv(opcode_type, 16#0A#),
      648 => to_slv(opcode_type, 16#0B#),
      649 => to_slv(opcode_type, 16#06#),
      650 => to_slv(opcode_type, 16#09#),
      651 => to_slv(opcode_type, 16#11#),
      652 => to_slv(opcode_type, 16#0B#),
      653 => to_slv(opcode_type, 16#07#),
      654 => to_slv(opcode_type, 16#11#),
      655 => to_slv(opcode_type, 16#0B#),
      656 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#02#),
      673 => to_slv(opcode_type, 16#09#),
      674 => to_slv(opcode_type, 16#09#),
      675 => to_slv(opcode_type, 16#06#),
      676 => to_slv(opcode_type, 16#0C#),
      677 => to_slv(opcode_type, 16#10#),
      678 => to_slv(opcode_type, 16#06#),
      679 => to_slv(opcode_type, 16#10#),
      680 => to_slv(opcode_type, 16#0D#),
      681 => to_slv(opcode_type, 16#06#),
      682 => to_slv(opcode_type, 16#07#),
      683 => to_slv(opcode_type, 16#0F#),
      684 => to_slv(opcode_type, 16#0E#),
      685 => to_slv(opcode_type, 16#06#),
      686 => to_slv(opcode_type, 16#0D#),
      687 => to_slv(opcode_type, 16#0D#),
      688 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#06#),
      705 => to_slv(opcode_type, 16#01#),
      706 => to_slv(opcode_type, 16#06#),
      707 => to_slv(opcode_type, 16#09#),
      708 => to_slv(opcode_type, 16#0D#),
      709 => to_slv(opcode_type, 16#0D#),
      710 => to_slv(opcode_type, 16#08#),
      711 => to_slv(opcode_type, 16#10#),
      712 => to_slv(opcode_type, 16#64#),
      713 => to_slv(opcode_type, 16#09#),
      714 => to_slv(opcode_type, 16#07#),
      715 => to_slv(opcode_type, 16#03#),
      716 => to_slv(opcode_type, 16#11#),
      717 => to_slv(opcode_type, 16#01#),
      718 => to_slv(opcode_type, 16#10#),
      719 => to_slv(opcode_type, 16#10#),
      720 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#01#),
      737 => to_slv(opcode_type, 16#07#),
      738 => to_slv(opcode_type, 16#08#),
      739 => to_slv(opcode_type, 16#09#),
      740 => to_slv(opcode_type, 16#10#),
      741 => to_slv(opcode_type, 16#0A#),
      742 => to_slv(opcode_type, 16#06#),
      743 => to_slv(opcode_type, 16#11#),
      744 => to_slv(opcode_type, 16#10#),
      745 => to_slv(opcode_type, 16#06#),
      746 => to_slv(opcode_type, 16#08#),
      747 => to_slv(opcode_type, 16#10#),
      748 => to_slv(opcode_type, 16#7E#),
      749 => to_slv(opcode_type, 16#08#),
      750 => to_slv(opcode_type, 16#7A#),
      751 => to_slv(opcode_type, 16#0B#),
      752 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#05#),
      769 => to_slv(opcode_type, 16#07#),
      770 => to_slv(opcode_type, 16#09#),
      771 => to_slv(opcode_type, 16#06#),
      772 => to_slv(opcode_type, 16#0A#),
      773 => to_slv(opcode_type, 16#0D#),
      774 => to_slv(opcode_type, 16#08#),
      775 => to_slv(opcode_type, 16#11#),
      776 => to_slv(opcode_type, 16#0F#),
      777 => to_slv(opcode_type, 16#06#),
      778 => to_slv(opcode_type, 16#08#),
      779 => to_slv(opcode_type, 16#10#),
      780 => to_slv(opcode_type, 16#0F#),
      781 => to_slv(opcode_type, 16#07#),
      782 => to_slv(opcode_type, 16#0F#),
      783 => to_slv(opcode_type, 16#0E#),
      784 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#03#),
      801 => to_slv(opcode_type, 16#08#),
      802 => to_slv(opcode_type, 16#09#),
      803 => to_slv(opcode_type, 16#07#),
      804 => to_slv(opcode_type, 16#15#),
      805 => to_slv(opcode_type, 16#0A#),
      806 => to_slv(opcode_type, 16#06#),
      807 => to_slv(opcode_type, 16#11#),
      808 => to_slv(opcode_type, 16#10#),
      809 => to_slv(opcode_type, 16#06#),
      810 => to_slv(opcode_type, 16#06#),
      811 => to_slv(opcode_type, 16#0B#),
      812 => to_slv(opcode_type, 16#0D#),
      813 => to_slv(opcode_type, 16#08#),
      814 => to_slv(opcode_type, 16#0C#),
      815 => to_slv(opcode_type, 16#0B#),
      816 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#09#),
      833 => to_slv(opcode_type, 16#02#),
      834 => to_slv(opcode_type, 16#07#),
      835 => to_slv(opcode_type, 16#04#),
      836 => to_slv(opcode_type, 16#10#),
      837 => to_slv(opcode_type, 16#03#),
      838 => to_slv(opcode_type, 16#0B#),
      839 => to_slv(opcode_type, 16#09#),
      840 => to_slv(opcode_type, 16#03#),
      841 => to_slv(opcode_type, 16#08#),
      842 => to_slv(opcode_type, 16#C6#),
      843 => to_slv(opcode_type, 16#0B#),
      844 => to_slv(opcode_type, 16#06#),
      845 => to_slv(opcode_type, 16#02#),
      846 => to_slv(opcode_type, 16#10#),
      847 => to_slv(opcode_type, 16#11#),
      848 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#04#),
      865 => to_slv(opcode_type, 16#08#),
      866 => to_slv(opcode_type, 16#08#),
      867 => to_slv(opcode_type, 16#09#),
      868 => to_slv(opcode_type, 16#0A#),
      869 => to_slv(opcode_type, 16#0C#),
      870 => to_slv(opcode_type, 16#09#),
      871 => to_slv(opcode_type, 16#0D#),
      872 => to_slv(opcode_type, 16#10#),
      873 => to_slv(opcode_type, 16#08#),
      874 => to_slv(opcode_type, 16#06#),
      875 => to_slv(opcode_type, 16#82#),
      876 => to_slv(opcode_type, 16#11#),
      877 => to_slv(opcode_type, 16#08#),
      878 => to_slv(opcode_type, 16#10#),
      879 => to_slv(opcode_type, 16#0C#),
      880 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#06#),
      897 => to_slv(opcode_type, 16#08#),
      898 => to_slv(opcode_type, 16#01#),
      899 => to_slv(opcode_type, 16#08#),
      900 => to_slv(opcode_type, 16#10#),
      901 => to_slv(opcode_type, 16#10#),
      902 => to_slv(opcode_type, 16#01#),
      903 => to_slv(opcode_type, 16#06#),
      904 => to_slv(opcode_type, 16#0D#),
      905 => to_slv(opcode_type, 16#0F#),
      906 => to_slv(opcode_type, 16#06#),
      907 => to_slv(opcode_type, 16#09#),
      908 => to_slv(opcode_type, 16#05#),
      909 => to_slv(opcode_type, 16#5B#),
      910 => to_slv(opcode_type, 16#0F#),
      911 => to_slv(opcode_type, 16#0F#),
      912 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#02#),
      929 => to_slv(opcode_type, 16#07#),
      930 => to_slv(opcode_type, 16#09#),
      931 => to_slv(opcode_type, 16#09#),
      932 => to_slv(opcode_type, 16#11#),
      933 => to_slv(opcode_type, 16#0E#),
      934 => to_slv(opcode_type, 16#07#),
      935 => to_slv(opcode_type, 16#0B#),
      936 => to_slv(opcode_type, 16#11#),
      937 => to_slv(opcode_type, 16#06#),
      938 => to_slv(opcode_type, 16#09#),
      939 => to_slv(opcode_type, 16#11#),
      940 => to_slv(opcode_type, 16#0C#),
      941 => to_slv(opcode_type, 16#08#),
      942 => to_slv(opcode_type, 16#0A#),
      943 => to_slv(opcode_type, 16#0A#),
      944 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#01#),
      961 => to_slv(opcode_type, 16#06#),
      962 => to_slv(opcode_type, 16#07#),
      963 => to_slv(opcode_type, 16#09#),
      964 => to_slv(opcode_type, 16#0E#),
      965 => to_slv(opcode_type, 16#0F#),
      966 => to_slv(opcode_type, 16#07#),
      967 => to_slv(opcode_type, 16#0F#),
      968 => to_slv(opcode_type, 16#0A#),
      969 => to_slv(opcode_type, 16#08#),
      970 => to_slv(opcode_type, 16#06#),
      971 => to_slv(opcode_type, 16#0D#),
      972 => to_slv(opcode_type, 16#11#),
      973 => to_slv(opcode_type, 16#09#),
      974 => to_slv(opcode_type, 16#0D#),
      975 => to_slv(opcode_type, 16#10#),
      976 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#02#),
      993 => to_slv(opcode_type, 16#08#),
      994 => to_slv(opcode_type, 16#08#),
      995 => to_slv(opcode_type, 16#06#),
      996 => to_slv(opcode_type, 16#10#),
      997 => to_slv(opcode_type, 16#10#),
      998 => to_slv(opcode_type, 16#06#),
      999 => to_slv(opcode_type, 16#0F#),
      1000 => to_slv(opcode_type, 16#0D#),
      1001 => to_slv(opcode_type, 16#06#),
      1002 => to_slv(opcode_type, 16#09#),
      1003 => to_slv(opcode_type, 16#0F#),
      1004 => to_slv(opcode_type, 16#10#),
      1005 => to_slv(opcode_type, 16#07#),
      1006 => to_slv(opcode_type, 16#0D#),
      1007 => to_slv(opcode_type, 16#0A#),
      1008 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#01#),
      1025 => to_slv(opcode_type, 16#08#),
      1026 => to_slv(opcode_type, 16#09#),
      1027 => to_slv(opcode_type, 16#06#),
      1028 => to_slv(opcode_type, 16#0E#),
      1029 => to_slv(opcode_type, 16#10#),
      1030 => to_slv(opcode_type, 16#06#),
      1031 => to_slv(opcode_type, 16#11#),
      1032 => to_slv(opcode_type, 16#0F#),
      1033 => to_slv(opcode_type, 16#09#),
      1034 => to_slv(opcode_type, 16#09#),
      1035 => to_slv(opcode_type, 16#0B#),
      1036 => to_slv(opcode_type, 16#0B#),
      1037 => to_slv(opcode_type, 16#08#),
      1038 => to_slv(opcode_type, 16#0D#),
      1039 => to_slv(opcode_type, 16#DF#),
      1040 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#09#),
      1057 => to_slv(opcode_type, 16#09#),
      1058 => to_slv(opcode_type, 16#06#),
      1059 => to_slv(opcode_type, 16#08#),
      1060 => to_slv(opcode_type, 16#0A#),
      1061 => to_slv(opcode_type, 16#10#),
      1062 => to_slv(opcode_type, 16#01#),
      1063 => to_slv(opcode_type, 16#0B#),
      1064 => to_slv(opcode_type, 16#01#),
      1065 => to_slv(opcode_type, 16#09#),
      1066 => to_slv(opcode_type, 16#0A#),
      1067 => to_slv(opcode_type, 16#0E#),
      1068 => to_slv(opcode_type, 16#03#),
      1069 => to_slv(opcode_type, 16#06#),
      1070 => to_slv(opcode_type, 16#10#),
      1071 => to_slv(opcode_type, 16#0F#),
      1072 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#09#),
      1089 => to_slv(opcode_type, 16#01#),
      1090 => to_slv(opcode_type, 16#01#),
      1091 => to_slv(opcode_type, 16#02#),
      1092 => to_slv(opcode_type, 16#0D#),
      1093 => to_slv(opcode_type, 16#06#),
      1094 => to_slv(opcode_type, 16#07#),
      1095 => to_slv(opcode_type, 16#04#),
      1096 => to_slv(opcode_type, 16#0E#),
      1097 => to_slv(opcode_type, 16#05#),
      1098 => to_slv(opcode_type, 16#0B#),
      1099 => to_slv(opcode_type, 16#09#),
      1100 => to_slv(opcode_type, 16#09#),
      1101 => to_slv(opcode_type, 16#0D#),
      1102 => to_slv(opcode_type, 16#0B#),
      1103 => to_slv(opcode_type, 16#0F#),
      1104 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#01#),
      1121 => to_slv(opcode_type, 16#08#),
      1122 => to_slv(opcode_type, 16#07#),
      1123 => to_slv(opcode_type, 16#08#),
      1124 => to_slv(opcode_type, 16#10#),
      1125 => to_slv(opcode_type, 16#11#),
      1126 => to_slv(opcode_type, 16#09#),
      1127 => to_slv(opcode_type, 16#0F#),
      1128 => to_slv(opcode_type, 16#11#),
      1129 => to_slv(opcode_type, 16#07#),
      1130 => to_slv(opcode_type, 16#08#),
      1131 => to_slv(opcode_type, 16#0A#),
      1132 => to_slv(opcode_type, 16#11#),
      1133 => to_slv(opcode_type, 16#09#),
      1134 => to_slv(opcode_type, 16#0F#),
      1135 => to_slv(opcode_type, 16#6D#),
      1136 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#07#),
      1153 => to_slv(opcode_type, 16#09#),
      1154 => to_slv(opcode_type, 16#01#),
      1155 => to_slv(opcode_type, 16#01#),
      1156 => to_slv(opcode_type, 16#0A#),
      1157 => to_slv(opcode_type, 16#08#),
      1158 => to_slv(opcode_type, 16#09#),
      1159 => to_slv(opcode_type, 16#10#),
      1160 => to_slv(opcode_type, 16#0C#),
      1161 => to_slv(opcode_type, 16#04#),
      1162 => to_slv(opcode_type, 16#11#),
      1163 => to_slv(opcode_type, 16#09#),
      1164 => to_slv(opcode_type, 16#07#),
      1165 => to_slv(opcode_type, 16#10#),
      1166 => to_slv(opcode_type, 16#0D#),
      1167 => to_slv(opcode_type, 16#32#),
      1168 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#07#),
      1185 => to_slv(opcode_type, 16#01#),
      1186 => to_slv(opcode_type, 16#03#),
      1187 => to_slv(opcode_type, 16#07#),
      1188 => to_slv(opcode_type, 16#10#),
      1189 => to_slv(opcode_type, 16#53#),
      1190 => to_slv(opcode_type, 16#07#),
      1191 => to_slv(opcode_type, 16#02#),
      1192 => to_slv(opcode_type, 16#06#),
      1193 => to_slv(opcode_type, 16#0D#),
      1194 => to_slv(opcode_type, 16#0B#),
      1195 => to_slv(opcode_type, 16#09#),
      1196 => to_slv(opcode_type, 16#02#),
      1197 => to_slv(opcode_type, 16#0A#),
      1198 => to_slv(opcode_type, 16#03#),
      1199 => to_slv(opcode_type, 16#0C#),
      1200 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#03#),
      1217 => to_slv(opcode_type, 16#07#),
      1218 => to_slv(opcode_type, 16#08#),
      1219 => to_slv(opcode_type, 16#06#),
      1220 => to_slv(opcode_type, 16#0D#),
      1221 => to_slv(opcode_type, 16#0F#),
      1222 => to_slv(opcode_type, 16#08#),
      1223 => to_slv(opcode_type, 16#10#),
      1224 => to_slv(opcode_type, 16#0A#),
      1225 => to_slv(opcode_type, 16#08#),
      1226 => to_slv(opcode_type, 16#09#),
      1227 => to_slv(opcode_type, 16#0E#),
      1228 => to_slv(opcode_type, 16#0A#),
      1229 => to_slv(opcode_type, 16#09#),
      1230 => to_slv(opcode_type, 16#0E#),
      1231 => to_slv(opcode_type, 16#0B#),
      1232 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#01#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#06#),
      1251 => to_slv(opcode_type, 16#07#),
      1252 => to_slv(opcode_type, 16#0E#),
      1253 => to_slv(opcode_type, 16#0C#),
      1254 => to_slv(opcode_type, 16#07#),
      1255 => to_slv(opcode_type, 16#0F#),
      1256 => to_slv(opcode_type, 16#0E#),
      1257 => to_slv(opcode_type, 16#08#),
      1258 => to_slv(opcode_type, 16#08#),
      1259 => to_slv(opcode_type, 16#0E#),
      1260 => to_slv(opcode_type, 16#0B#),
      1261 => to_slv(opcode_type, 16#08#),
      1262 => to_slv(opcode_type, 16#0F#),
      1263 => to_slv(opcode_type, 16#70#),
      1264 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#04#),
      1281 => to_slv(opcode_type, 16#07#),
      1282 => to_slv(opcode_type, 16#07#),
      1283 => to_slv(opcode_type, 16#06#),
      1284 => to_slv(opcode_type, 16#0A#),
      1285 => to_slv(opcode_type, 16#10#),
      1286 => to_slv(opcode_type, 16#08#),
      1287 => to_slv(opcode_type, 16#0B#),
      1288 => to_slv(opcode_type, 16#0B#),
      1289 => to_slv(opcode_type, 16#07#),
      1290 => to_slv(opcode_type, 16#08#),
      1291 => to_slv(opcode_type, 16#0F#),
      1292 => to_slv(opcode_type, 16#0B#),
      1293 => to_slv(opcode_type, 16#07#),
      1294 => to_slv(opcode_type, 16#0E#),
      1295 => to_slv(opcode_type, 16#0B#),
      1296 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#05#),
      1313 => to_slv(opcode_type, 16#07#),
      1314 => to_slv(opcode_type, 16#09#),
      1315 => to_slv(opcode_type, 16#08#),
      1316 => to_slv(opcode_type, 16#0C#),
      1317 => to_slv(opcode_type, 16#EB#),
      1318 => to_slv(opcode_type, 16#06#),
      1319 => to_slv(opcode_type, 16#0D#),
      1320 => to_slv(opcode_type, 16#0E#),
      1321 => to_slv(opcode_type, 16#06#),
      1322 => to_slv(opcode_type, 16#09#),
      1323 => to_slv(opcode_type, 16#0F#),
      1324 => to_slv(opcode_type, 16#0E#),
      1325 => to_slv(opcode_type, 16#06#),
      1326 => to_slv(opcode_type, 16#0E#),
      1327 => to_slv(opcode_type, 16#0E#),
      1328 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#06#),
      1345 => to_slv(opcode_type, 16#07#),
      1346 => to_slv(opcode_type, 16#06#),
      1347 => to_slv(opcode_type, 16#04#),
      1348 => to_slv(opcode_type, 16#0B#),
      1349 => to_slv(opcode_type, 16#03#),
      1350 => to_slv(opcode_type, 16#11#),
      1351 => to_slv(opcode_type, 16#08#),
      1352 => to_slv(opcode_type, 16#09#),
      1353 => to_slv(opcode_type, 16#10#),
      1354 => to_slv(opcode_type, 16#0F#),
      1355 => to_slv(opcode_type, 16#02#),
      1356 => to_slv(opcode_type, 16#0E#),
      1357 => to_slv(opcode_type, 16#02#),
      1358 => to_slv(opcode_type, 16#05#),
      1359 => to_slv(opcode_type, 16#0D#),
      1360 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#02#),
      1377 => to_slv(opcode_type, 16#08#),
      1378 => to_slv(opcode_type, 16#06#),
      1379 => to_slv(opcode_type, 16#06#),
      1380 => to_slv(opcode_type, 16#0D#),
      1381 => to_slv(opcode_type, 16#0B#),
      1382 => to_slv(opcode_type, 16#08#),
      1383 => to_slv(opcode_type, 16#11#),
      1384 => to_slv(opcode_type, 16#11#),
      1385 => to_slv(opcode_type, 16#08#),
      1386 => to_slv(opcode_type, 16#09#),
      1387 => to_slv(opcode_type, 16#54#),
      1388 => to_slv(opcode_type, 16#0C#),
      1389 => to_slv(opcode_type, 16#06#),
      1390 => to_slv(opcode_type, 16#81#),
      1391 => to_slv(opcode_type, 16#10#),
      1392 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#05#),
      1409 => to_slv(opcode_type, 16#07#),
      1410 => to_slv(opcode_type, 16#07#),
      1411 => to_slv(opcode_type, 16#09#),
      1412 => to_slv(opcode_type, 16#DD#),
      1413 => to_slv(opcode_type, 16#0B#),
      1414 => to_slv(opcode_type, 16#08#),
      1415 => to_slv(opcode_type, 16#0A#),
      1416 => to_slv(opcode_type, 16#11#),
      1417 => to_slv(opcode_type, 16#08#),
      1418 => to_slv(opcode_type, 16#08#),
      1419 => to_slv(opcode_type, 16#11#),
      1420 => to_slv(opcode_type, 16#0A#),
      1421 => to_slv(opcode_type, 16#09#),
      1422 => to_slv(opcode_type, 16#11#),
      1423 => to_slv(opcode_type, 16#0D#),
      1424 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#08#),
      1441 => to_slv(opcode_type, 16#03#),
      1442 => to_slv(opcode_type, 16#04#),
      1443 => to_slv(opcode_type, 16#09#),
      1444 => to_slv(opcode_type, 16#0E#),
      1445 => to_slv(opcode_type, 16#0A#),
      1446 => to_slv(opcode_type, 16#06#),
      1447 => to_slv(opcode_type, 16#06#),
      1448 => to_slv(opcode_type, 16#05#),
      1449 => to_slv(opcode_type, 16#10#),
      1450 => to_slv(opcode_type, 16#09#),
      1451 => to_slv(opcode_type, 16#0D#),
      1452 => to_slv(opcode_type, 16#0F#),
      1453 => to_slv(opcode_type, 16#04#),
      1454 => to_slv(opcode_type, 16#05#),
      1455 => to_slv(opcode_type, 16#11#),
      1456 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#05#),
      1473 => to_slv(opcode_type, 16#07#),
      1474 => to_slv(opcode_type, 16#06#),
      1475 => to_slv(opcode_type, 16#06#),
      1476 => to_slv(opcode_type, 16#0C#),
      1477 => to_slv(opcode_type, 16#0B#),
      1478 => to_slv(opcode_type, 16#07#),
      1479 => to_slv(opcode_type, 16#11#),
      1480 => to_slv(opcode_type, 16#10#),
      1481 => to_slv(opcode_type, 16#08#),
      1482 => to_slv(opcode_type, 16#06#),
      1483 => to_slv(opcode_type, 16#11#),
      1484 => to_slv(opcode_type, 16#10#),
      1485 => to_slv(opcode_type, 16#07#),
      1486 => to_slv(opcode_type, 16#87#),
      1487 => to_slv(opcode_type, 16#0F#),
      1488 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#03#),
      1505 => to_slv(opcode_type, 16#08#),
      1506 => to_slv(opcode_type, 16#08#),
      1507 => to_slv(opcode_type, 16#08#),
      1508 => to_slv(opcode_type, 16#0D#),
      1509 => to_slv(opcode_type, 16#0A#),
      1510 => to_slv(opcode_type, 16#06#),
      1511 => to_slv(opcode_type, 16#0A#),
      1512 => to_slv(opcode_type, 16#0E#),
      1513 => to_slv(opcode_type, 16#06#),
      1514 => to_slv(opcode_type, 16#08#),
      1515 => to_slv(opcode_type, 16#0D#),
      1516 => to_slv(opcode_type, 16#0C#),
      1517 => to_slv(opcode_type, 16#08#),
      1518 => to_slv(opcode_type, 16#0A#),
      1519 => to_slv(opcode_type, 16#0C#),
      1520 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#06#),
      1537 => to_slv(opcode_type, 16#01#),
      1538 => to_slv(opcode_type, 16#05#),
      1539 => to_slv(opcode_type, 16#04#),
      1540 => to_slv(opcode_type, 16#11#),
      1541 => to_slv(opcode_type, 16#08#),
      1542 => to_slv(opcode_type, 16#06#),
      1543 => to_slv(opcode_type, 16#01#),
      1544 => to_slv(opcode_type, 16#0D#),
      1545 => to_slv(opcode_type, 16#04#),
      1546 => to_slv(opcode_type, 16#0B#),
      1547 => to_slv(opcode_type, 16#06#),
      1548 => to_slv(opcode_type, 16#04#),
      1549 => to_slv(opcode_type, 16#0F#),
      1550 => to_slv(opcode_type, 16#04#),
      1551 => to_slv(opcode_type, 16#11#),
      1552 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#04#),
      1569 => to_slv(opcode_type, 16#09#),
      1570 => to_slv(opcode_type, 16#08#),
      1571 => to_slv(opcode_type, 16#09#),
      1572 => to_slv(opcode_type, 16#11#),
      1573 => to_slv(opcode_type, 16#0B#),
      1574 => to_slv(opcode_type, 16#06#),
      1575 => to_slv(opcode_type, 16#0F#),
      1576 => to_slv(opcode_type, 16#0B#),
      1577 => to_slv(opcode_type, 16#09#),
      1578 => to_slv(opcode_type, 16#08#),
      1579 => to_slv(opcode_type, 16#0E#),
      1580 => to_slv(opcode_type, 16#0A#),
      1581 => to_slv(opcode_type, 16#06#),
      1582 => to_slv(opcode_type, 16#11#),
      1583 => to_slv(opcode_type, 16#0D#),
      1584 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#09#),
      1601 => to_slv(opcode_type, 16#02#),
      1602 => to_slv(opcode_type, 16#05#),
      1603 => to_slv(opcode_type, 16#06#),
      1604 => to_slv(opcode_type, 16#0F#),
      1605 => to_slv(opcode_type, 16#0B#),
      1606 => to_slv(opcode_type, 16#08#),
      1607 => to_slv(opcode_type, 16#03#),
      1608 => to_slv(opcode_type, 16#08#),
      1609 => to_slv(opcode_type, 16#0C#),
      1610 => to_slv(opcode_type, 16#0C#),
      1611 => to_slv(opcode_type, 16#08#),
      1612 => to_slv(opcode_type, 16#07#),
      1613 => to_slv(opcode_type, 16#51#),
      1614 => to_slv(opcode_type, 16#10#),
      1615 => to_slv(opcode_type, 16#0A#),
      1616 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#09#),
      1633 => to_slv(opcode_type, 16#01#),
      1634 => to_slv(opcode_type, 16#06#),
      1635 => to_slv(opcode_type, 16#04#),
      1636 => to_slv(opcode_type, 16#11#),
      1637 => to_slv(opcode_type, 16#03#),
      1638 => to_slv(opcode_type, 16#10#),
      1639 => to_slv(opcode_type, 16#09#),
      1640 => to_slv(opcode_type, 16#01#),
      1641 => to_slv(opcode_type, 16#03#),
      1642 => to_slv(opcode_type, 16#0A#),
      1643 => to_slv(opcode_type, 16#06#),
      1644 => to_slv(opcode_type, 16#07#),
      1645 => to_slv(opcode_type, 16#11#),
      1646 => to_slv(opcode_type, 16#0F#),
      1647 => to_slv(opcode_type, 16#0B#),
      1648 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#01#),
      1666 => to_slv(opcode_type, 16#02#),
      1667 => to_slv(opcode_type, 16#01#),
      1668 => to_slv(opcode_type, 16#0C#),
      1669 => to_slv(opcode_type, 16#06#),
      1670 => to_slv(opcode_type, 16#05#),
      1671 => to_slv(opcode_type, 16#06#),
      1672 => to_slv(opcode_type, 16#0E#),
      1673 => to_slv(opcode_type, 16#0C#),
      1674 => to_slv(opcode_type, 16#07#),
      1675 => to_slv(opcode_type, 16#08#),
      1676 => to_slv(opcode_type, 16#0A#),
      1677 => to_slv(opcode_type, 16#11#),
      1678 => to_slv(opcode_type, 16#04#),
      1679 => to_slv(opcode_type, 16#0A#),
      1680 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#05#),
      1697 => to_slv(opcode_type, 16#08#),
      1698 => to_slv(opcode_type, 16#09#),
      1699 => to_slv(opcode_type, 16#07#),
      1700 => to_slv(opcode_type, 16#0B#),
      1701 => to_slv(opcode_type, 16#10#),
      1702 => to_slv(opcode_type, 16#07#),
      1703 => to_slv(opcode_type, 16#0F#),
      1704 => to_slv(opcode_type, 16#0C#),
      1705 => to_slv(opcode_type, 16#08#),
      1706 => to_slv(opcode_type, 16#06#),
      1707 => to_slv(opcode_type, 16#0D#),
      1708 => to_slv(opcode_type, 16#0C#),
      1709 => to_slv(opcode_type, 16#06#),
      1710 => to_slv(opcode_type, 16#11#),
      1711 => to_slv(opcode_type, 16#10#),
      1712 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#04#),
      1729 => to_slv(opcode_type, 16#07#),
      1730 => to_slv(opcode_type, 16#06#),
      1731 => to_slv(opcode_type, 16#09#),
      1732 => to_slv(opcode_type, 16#10#),
      1733 => to_slv(opcode_type, 16#0E#),
      1734 => to_slv(opcode_type, 16#09#),
      1735 => to_slv(opcode_type, 16#11#),
      1736 => to_slv(opcode_type, 16#0A#),
      1737 => to_slv(opcode_type, 16#09#),
      1738 => to_slv(opcode_type, 16#08#),
      1739 => to_slv(opcode_type, 16#0F#),
      1740 => to_slv(opcode_type, 16#0A#),
      1741 => to_slv(opcode_type, 16#08#),
      1742 => to_slv(opcode_type, 16#11#),
      1743 => to_slv(opcode_type, 16#0C#),
      1744 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#09#),
      1761 => to_slv(opcode_type, 16#05#),
      1762 => to_slv(opcode_type, 16#03#),
      1763 => to_slv(opcode_type, 16#07#),
      1764 => to_slv(opcode_type, 16#0F#),
      1765 => to_slv(opcode_type, 16#0F#),
      1766 => to_slv(opcode_type, 16#08#),
      1767 => to_slv(opcode_type, 16#09#),
      1768 => to_slv(opcode_type, 16#06#),
      1769 => to_slv(opcode_type, 16#0F#),
      1770 => to_slv(opcode_type, 16#0F#),
      1771 => to_slv(opcode_type, 16#04#),
      1772 => to_slv(opcode_type, 16#0F#),
      1773 => to_slv(opcode_type, 16#01#),
      1774 => to_slv(opcode_type, 16#03#),
      1775 => to_slv(opcode_type, 16#0B#),
      1776 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#01#),
      1793 => to_slv(opcode_type, 16#07#),
      1794 => to_slv(opcode_type, 16#06#),
      1795 => to_slv(opcode_type, 16#09#),
      1796 => to_slv(opcode_type, 16#10#),
      1797 => to_slv(opcode_type, 16#0C#),
      1798 => to_slv(opcode_type, 16#08#),
      1799 => to_slv(opcode_type, 16#10#),
      1800 => to_slv(opcode_type, 16#0C#),
      1801 => to_slv(opcode_type, 16#06#),
      1802 => to_slv(opcode_type, 16#09#),
      1803 => to_slv(opcode_type, 16#0A#),
      1804 => to_slv(opcode_type, 16#0C#),
      1805 => to_slv(opcode_type, 16#06#),
      1806 => to_slv(opcode_type, 16#0D#),
      1807 => to_slv(opcode_type, 16#0D#),
      1808 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#06#),
      1825 => to_slv(opcode_type, 16#07#),
      1826 => to_slv(opcode_type, 16#05#),
      1827 => to_slv(opcode_type, 16#09#),
      1828 => to_slv(opcode_type, 16#0C#),
      1829 => to_slv(opcode_type, 16#10#),
      1830 => to_slv(opcode_type, 16#04#),
      1831 => to_slv(opcode_type, 16#04#),
      1832 => to_slv(opcode_type, 16#11#),
      1833 => to_slv(opcode_type, 16#07#),
      1834 => to_slv(opcode_type, 16#07#),
      1835 => to_slv(opcode_type, 16#03#),
      1836 => to_slv(opcode_type, 16#0B#),
      1837 => to_slv(opcode_type, 16#02#),
      1838 => to_slv(opcode_type, 16#0F#),
      1839 => to_slv(opcode_type, 16#0B#),
      1840 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#01#),
      1857 => to_slv(opcode_type, 16#09#),
      1858 => to_slv(opcode_type, 16#09#),
      1859 => to_slv(opcode_type, 16#08#),
      1860 => to_slv(opcode_type, 16#10#),
      1861 => to_slv(opcode_type, 16#10#),
      1862 => to_slv(opcode_type, 16#06#),
      1863 => to_slv(opcode_type, 16#10#),
      1864 => to_slv(opcode_type, 16#0F#),
      1865 => to_slv(opcode_type, 16#06#),
      1866 => to_slv(opcode_type, 16#08#),
      1867 => to_slv(opcode_type, 16#0B#),
      1868 => to_slv(opcode_type, 16#0C#),
      1869 => to_slv(opcode_type, 16#07#),
      1870 => to_slv(opcode_type, 16#0E#),
      1871 => to_slv(opcode_type, 16#11#),
      1872 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#02#),
      1889 => to_slv(opcode_type, 16#08#),
      1890 => to_slv(opcode_type, 16#09#),
      1891 => to_slv(opcode_type, 16#09#),
      1892 => to_slv(opcode_type, 16#0D#),
      1893 => to_slv(opcode_type, 16#0A#),
      1894 => to_slv(opcode_type, 16#09#),
      1895 => to_slv(opcode_type, 16#0B#),
      1896 => to_slv(opcode_type, 16#0C#),
      1897 => to_slv(opcode_type, 16#09#),
      1898 => to_slv(opcode_type, 16#08#),
      1899 => to_slv(opcode_type, 16#0B#),
      1900 => to_slv(opcode_type, 16#B7#),
      1901 => to_slv(opcode_type, 16#08#),
      1902 => to_slv(opcode_type, 16#0F#),
      1903 => to_slv(opcode_type, 16#11#),
      1904 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#03#),
      1921 => to_slv(opcode_type, 16#08#),
      1922 => to_slv(opcode_type, 16#08#),
      1923 => to_slv(opcode_type, 16#08#),
      1924 => to_slv(opcode_type, 16#10#),
      1925 => to_slv(opcode_type, 16#0A#),
      1926 => to_slv(opcode_type, 16#09#),
      1927 => to_slv(opcode_type, 16#0B#),
      1928 => to_slv(opcode_type, 16#0A#),
      1929 => to_slv(opcode_type, 16#09#),
      1930 => to_slv(opcode_type, 16#07#),
      1931 => to_slv(opcode_type, 16#61#),
      1932 => to_slv(opcode_type, 16#24#),
      1933 => to_slv(opcode_type, 16#06#),
      1934 => to_slv(opcode_type, 16#0F#),
      1935 => to_slv(opcode_type, 16#D2#),
      1936 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#01#),
      1953 => to_slv(opcode_type, 16#08#),
      1954 => to_slv(opcode_type, 16#07#),
      1955 => to_slv(opcode_type, 16#07#),
      1956 => to_slv(opcode_type, 16#0D#),
      1957 => to_slv(opcode_type, 16#0C#),
      1958 => to_slv(opcode_type, 16#07#),
      1959 => to_slv(opcode_type, 16#0F#),
      1960 => to_slv(opcode_type, 16#0F#),
      1961 => to_slv(opcode_type, 16#06#),
      1962 => to_slv(opcode_type, 16#06#),
      1963 => to_slv(opcode_type, 16#0C#),
      1964 => to_slv(opcode_type, 16#0F#),
      1965 => to_slv(opcode_type, 16#09#),
      1966 => to_slv(opcode_type, 16#60#),
      1967 => to_slv(opcode_type, 16#0B#),
      1968 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#06#),
      1985 => to_slv(opcode_type, 16#08#),
      1986 => to_slv(opcode_type, 16#08#),
      1987 => to_slv(opcode_type, 16#02#),
      1988 => to_slv(opcode_type, 16#0D#),
      1989 => to_slv(opcode_type, 16#07#),
      1990 => to_slv(opcode_type, 16#0B#),
      1991 => to_slv(opcode_type, 16#93#),
      1992 => to_slv(opcode_type, 16#04#),
      1993 => to_slv(opcode_type, 16#09#),
      1994 => to_slv(opcode_type, 16#0E#),
      1995 => to_slv(opcode_type, 16#71#),
      1996 => to_slv(opcode_type, 16#06#),
      1997 => to_slv(opcode_type, 16#03#),
      1998 => to_slv(opcode_type, 16#0B#),
      1999 => to_slv(opcode_type, 16#B3#),
      2000 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#05#),
      2017 => to_slv(opcode_type, 16#08#),
      2018 => to_slv(opcode_type, 16#09#),
      2019 => to_slv(opcode_type, 16#08#),
      2020 => to_slv(opcode_type, 16#0D#),
      2021 => to_slv(opcode_type, 16#6D#),
      2022 => to_slv(opcode_type, 16#08#),
      2023 => to_slv(opcode_type, 16#0E#),
      2024 => to_slv(opcode_type, 16#0A#),
      2025 => to_slv(opcode_type, 16#06#),
      2026 => to_slv(opcode_type, 16#08#),
      2027 => to_slv(opcode_type, 16#10#),
      2028 => to_slv(opcode_type, 16#11#),
      2029 => to_slv(opcode_type, 16#06#),
      2030 => to_slv(opcode_type, 16#0F#),
      2031 => to_slv(opcode_type, 16#0F#),
      2032 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#01#),
      2049 => to_slv(opcode_type, 16#06#),
      2050 => to_slv(opcode_type, 16#07#),
      2051 => to_slv(opcode_type, 16#07#),
      2052 => to_slv(opcode_type, 16#0A#),
      2053 => to_slv(opcode_type, 16#11#),
      2054 => to_slv(opcode_type, 16#07#),
      2055 => to_slv(opcode_type, 16#0D#),
      2056 => to_slv(opcode_type, 16#11#),
      2057 => to_slv(opcode_type, 16#06#),
      2058 => to_slv(opcode_type, 16#09#),
      2059 => to_slv(opcode_type, 16#10#),
      2060 => to_slv(opcode_type, 16#2F#),
      2061 => to_slv(opcode_type, 16#07#),
      2062 => to_slv(opcode_type, 16#25#),
      2063 => to_slv(opcode_type, 16#0C#),
      2064 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#09#),
      2081 => to_slv(opcode_type, 16#05#),
      2082 => to_slv(opcode_type, 16#09#),
      2083 => to_slv(opcode_type, 16#07#),
      2084 => to_slv(opcode_type, 16#0C#),
      2085 => to_slv(opcode_type, 16#0D#),
      2086 => to_slv(opcode_type, 16#06#),
      2087 => to_slv(opcode_type, 16#16#),
      2088 => to_slv(opcode_type, 16#0A#),
      2089 => to_slv(opcode_type, 16#09#),
      2090 => to_slv(opcode_type, 16#07#),
      2091 => to_slv(opcode_type, 16#06#),
      2092 => to_slv(opcode_type, 16#10#),
      2093 => to_slv(opcode_type, 16#0E#),
      2094 => to_slv(opcode_type, 16#11#),
      2095 => to_slv(opcode_type, 16#43#),
      2096 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#03#),
      2113 => to_slv(opcode_type, 16#07#),
      2114 => to_slv(opcode_type, 16#09#),
      2115 => to_slv(opcode_type, 16#07#),
      2116 => to_slv(opcode_type, 16#0F#),
      2117 => to_slv(opcode_type, 16#11#),
      2118 => to_slv(opcode_type, 16#06#),
      2119 => to_slv(opcode_type, 16#10#),
      2120 => to_slv(opcode_type, 16#A9#),
      2121 => to_slv(opcode_type, 16#08#),
      2122 => to_slv(opcode_type, 16#08#),
      2123 => to_slv(opcode_type, 16#0F#),
      2124 => to_slv(opcode_type, 16#0D#),
      2125 => to_slv(opcode_type, 16#06#),
      2126 => to_slv(opcode_type, 16#0C#),
      2127 => to_slv(opcode_type, 16#0D#),
      2128 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#09#),
      2146 => to_slv(opcode_type, 16#05#),
      2147 => to_slv(opcode_type, 16#04#),
      2148 => to_slv(opcode_type, 16#0A#),
      2149 => to_slv(opcode_type, 16#04#),
      2150 => to_slv(opcode_type, 16#04#),
      2151 => to_slv(opcode_type, 16#10#),
      2152 => to_slv(opcode_type, 16#08#),
      2153 => to_slv(opcode_type, 16#04#),
      2154 => to_slv(opcode_type, 16#01#),
      2155 => to_slv(opcode_type, 16#0D#),
      2156 => to_slv(opcode_type, 16#08#),
      2157 => to_slv(opcode_type, 16#01#),
      2158 => to_slv(opcode_type, 16#3D#),
      2159 => to_slv(opcode_type, 16#0C#),
      2160 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#05#),
      2177 => to_slv(opcode_type, 16#07#),
      2178 => to_slv(opcode_type, 16#06#),
      2179 => to_slv(opcode_type, 16#07#),
      2180 => to_slv(opcode_type, 16#0A#),
      2181 => to_slv(opcode_type, 16#0F#),
      2182 => to_slv(opcode_type, 16#08#),
      2183 => to_slv(opcode_type, 16#10#),
      2184 => to_slv(opcode_type, 16#AE#),
      2185 => to_slv(opcode_type, 16#07#),
      2186 => to_slv(opcode_type, 16#09#),
      2187 => to_slv(opcode_type, 16#10#),
      2188 => to_slv(opcode_type, 16#0F#),
      2189 => to_slv(opcode_type, 16#09#),
      2190 => to_slv(opcode_type, 16#11#),
      2191 => to_slv(opcode_type, 16#0A#),
      2192 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#08#),
      2209 => to_slv(opcode_type, 16#06#),
      2210 => to_slv(opcode_type, 16#01#),
      2211 => to_slv(opcode_type, 16#07#),
      2212 => to_slv(opcode_type, 16#0A#),
      2213 => to_slv(opcode_type, 16#0C#),
      2214 => to_slv(opcode_type, 16#04#),
      2215 => to_slv(opcode_type, 16#08#),
      2216 => to_slv(opcode_type, 16#0C#),
      2217 => to_slv(opcode_type, 16#11#),
      2218 => to_slv(opcode_type, 16#06#),
      2219 => to_slv(opcode_type, 16#08#),
      2220 => to_slv(opcode_type, 16#04#),
      2221 => to_slv(opcode_type, 16#0E#),
      2222 => to_slv(opcode_type, 16#0E#),
      2223 => to_slv(opcode_type, 16#0D#),
      2224 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#03#),
      2241 => to_slv(opcode_type, 16#07#),
      2242 => to_slv(opcode_type, 16#06#),
      2243 => to_slv(opcode_type, 16#09#),
      2244 => to_slv(opcode_type, 16#0A#),
      2245 => to_slv(opcode_type, 16#0B#),
      2246 => to_slv(opcode_type, 16#08#),
      2247 => to_slv(opcode_type, 16#0F#),
      2248 => to_slv(opcode_type, 16#0F#),
      2249 => to_slv(opcode_type, 16#09#),
      2250 => to_slv(opcode_type, 16#07#),
      2251 => to_slv(opcode_type, 16#0B#),
      2252 => to_slv(opcode_type, 16#11#),
      2253 => to_slv(opcode_type, 16#07#),
      2254 => to_slv(opcode_type, 16#0C#),
      2255 => to_slv(opcode_type, 16#10#),
      2256 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#09#),
      2273 => to_slv(opcode_type, 16#05#),
      2274 => to_slv(opcode_type, 16#07#),
      2275 => to_slv(opcode_type, 16#07#),
      2276 => to_slv(opcode_type, 16#0F#),
      2277 => to_slv(opcode_type, 16#0C#),
      2278 => to_slv(opcode_type, 16#04#),
      2279 => to_slv(opcode_type, 16#11#),
      2280 => to_slv(opcode_type, 16#04#),
      2281 => to_slv(opcode_type, 16#07#),
      2282 => to_slv(opcode_type, 16#09#),
      2283 => to_slv(opcode_type, 16#0A#),
      2284 => to_slv(opcode_type, 16#9D#),
      2285 => to_slv(opcode_type, 16#06#),
      2286 => to_slv(opcode_type, 16#10#),
      2287 => to_slv(opcode_type, 16#0D#),
      2288 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#03#),
      2305 => to_slv(opcode_type, 16#07#),
      2306 => to_slv(opcode_type, 16#09#),
      2307 => to_slv(opcode_type, 16#06#),
      2308 => to_slv(opcode_type, 16#10#),
      2309 => to_slv(opcode_type, 16#0E#),
      2310 => to_slv(opcode_type, 16#06#),
      2311 => to_slv(opcode_type, 16#0C#),
      2312 => to_slv(opcode_type, 16#0F#),
      2313 => to_slv(opcode_type, 16#09#),
      2314 => to_slv(opcode_type, 16#07#),
      2315 => to_slv(opcode_type, 16#0E#),
      2316 => to_slv(opcode_type, 16#0C#),
      2317 => to_slv(opcode_type, 16#06#),
      2318 => to_slv(opcode_type, 16#0E#),
      2319 => to_slv(opcode_type, 16#11#),
      2320 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#04#),
      2337 => to_slv(opcode_type, 16#08#),
      2338 => to_slv(opcode_type, 16#08#),
      2339 => to_slv(opcode_type, 16#07#),
      2340 => to_slv(opcode_type, 16#0D#),
      2341 => to_slv(opcode_type, 16#0D#),
      2342 => to_slv(opcode_type, 16#08#),
      2343 => to_slv(opcode_type, 16#0A#),
      2344 => to_slv(opcode_type, 16#11#),
      2345 => to_slv(opcode_type, 16#08#),
      2346 => to_slv(opcode_type, 16#08#),
      2347 => to_slv(opcode_type, 16#11#),
      2348 => to_slv(opcode_type, 16#0F#),
      2349 => to_slv(opcode_type, 16#07#),
      2350 => to_slv(opcode_type, 16#10#),
      2351 => to_slv(opcode_type, 16#0B#),
      2352 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#01#),
      2369 => to_slv(opcode_type, 16#08#),
      2370 => to_slv(opcode_type, 16#09#),
      2371 => to_slv(opcode_type, 16#08#),
      2372 => to_slv(opcode_type, 16#0F#),
      2373 => to_slv(opcode_type, 16#0F#),
      2374 => to_slv(opcode_type, 16#06#),
      2375 => to_slv(opcode_type, 16#A6#),
      2376 => to_slv(opcode_type, 16#0E#),
      2377 => to_slv(opcode_type, 16#08#),
      2378 => to_slv(opcode_type, 16#09#),
      2379 => to_slv(opcode_type, 16#0D#),
      2380 => to_slv(opcode_type, 16#0A#),
      2381 => to_slv(opcode_type, 16#09#),
      2382 => to_slv(opcode_type, 16#10#),
      2383 => to_slv(opcode_type, 16#0C#),
      2384 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#01#),
      2401 => to_slv(opcode_type, 16#08#),
      2402 => to_slv(opcode_type, 16#09#),
      2403 => to_slv(opcode_type, 16#06#),
      2404 => to_slv(opcode_type, 16#11#),
      2405 => to_slv(opcode_type, 16#0E#),
      2406 => to_slv(opcode_type, 16#08#),
      2407 => to_slv(opcode_type, 16#0E#),
      2408 => to_slv(opcode_type, 16#0D#),
      2409 => to_slv(opcode_type, 16#09#),
      2410 => to_slv(opcode_type, 16#09#),
      2411 => to_slv(opcode_type, 16#E5#),
      2412 => to_slv(opcode_type, 16#AA#),
      2413 => to_slv(opcode_type, 16#07#),
      2414 => to_slv(opcode_type, 16#0C#),
      2415 => to_slv(opcode_type, 16#11#),
      2416 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#01#),
      2433 => to_slv(opcode_type, 16#09#),
      2434 => to_slv(opcode_type, 16#07#),
      2435 => to_slv(opcode_type, 16#06#),
      2436 => to_slv(opcode_type, 16#0F#),
      2437 => to_slv(opcode_type, 16#0A#),
      2438 => to_slv(opcode_type, 16#07#),
      2439 => to_slv(opcode_type, 16#0E#),
      2440 => to_slv(opcode_type, 16#10#),
      2441 => to_slv(opcode_type, 16#06#),
      2442 => to_slv(opcode_type, 16#09#),
      2443 => to_slv(opcode_type, 16#0F#),
      2444 => to_slv(opcode_type, 16#0F#),
      2445 => to_slv(opcode_type, 16#08#),
      2446 => to_slv(opcode_type, 16#EC#),
      2447 => to_slv(opcode_type, 16#0B#),
      2448 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#01#),
      2465 => to_slv(opcode_type, 16#06#),
      2466 => to_slv(opcode_type, 16#07#),
      2467 => to_slv(opcode_type, 16#06#),
      2468 => to_slv(opcode_type, 16#0A#),
      2469 => to_slv(opcode_type, 16#0A#),
      2470 => to_slv(opcode_type, 16#06#),
      2471 => to_slv(opcode_type, 16#0F#),
      2472 => to_slv(opcode_type, 16#11#),
      2473 => to_slv(opcode_type, 16#09#),
      2474 => to_slv(opcode_type, 16#09#),
      2475 => to_slv(opcode_type, 16#A6#),
      2476 => to_slv(opcode_type, 16#A8#),
      2477 => to_slv(opcode_type, 16#07#),
      2478 => to_slv(opcode_type, 16#0D#),
      2479 => to_slv(opcode_type, 16#0F#),
      2480 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#01#),
      2497 => to_slv(opcode_type, 16#06#),
      2498 => to_slv(opcode_type, 16#06#),
      2499 => to_slv(opcode_type, 16#07#),
      2500 => to_slv(opcode_type, 16#11#),
      2501 => to_slv(opcode_type, 16#0C#),
      2502 => to_slv(opcode_type, 16#07#),
      2503 => to_slv(opcode_type, 16#11#),
      2504 => to_slv(opcode_type, 16#0B#),
      2505 => to_slv(opcode_type, 16#09#),
      2506 => to_slv(opcode_type, 16#07#),
      2507 => to_slv(opcode_type, 16#10#),
      2508 => to_slv(opcode_type, 16#0A#),
      2509 => to_slv(opcode_type, 16#06#),
      2510 => to_slv(opcode_type, 16#10#),
      2511 => to_slv(opcode_type, 16#11#),
      2512 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#08#),
      2529 => to_slv(opcode_type, 16#02#),
      2530 => to_slv(opcode_type, 16#03#),
      2531 => to_slv(opcode_type, 16#05#),
      2532 => to_slv(opcode_type, 16#1E#),
      2533 => to_slv(opcode_type, 16#06#),
      2534 => to_slv(opcode_type, 16#01#),
      2535 => to_slv(opcode_type, 16#02#),
      2536 => to_slv(opcode_type, 16#0C#),
      2537 => to_slv(opcode_type, 16#08#),
      2538 => to_slv(opcode_type, 16#06#),
      2539 => to_slv(opcode_type, 16#0E#),
      2540 => to_slv(opcode_type, 16#0B#),
      2541 => to_slv(opcode_type, 16#06#),
      2542 => to_slv(opcode_type, 16#6C#),
      2543 => to_slv(opcode_type, 16#0F#),
      2544 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#03#),
      2561 => to_slv(opcode_type, 16#07#),
      2562 => to_slv(opcode_type, 16#06#),
      2563 => to_slv(opcode_type, 16#06#),
      2564 => to_slv(opcode_type, 16#F5#),
      2565 => to_slv(opcode_type, 16#11#),
      2566 => to_slv(opcode_type, 16#09#),
      2567 => to_slv(opcode_type, 16#11#),
      2568 => to_slv(opcode_type, 16#11#),
      2569 => to_slv(opcode_type, 16#09#),
      2570 => to_slv(opcode_type, 16#06#),
      2571 => to_slv(opcode_type, 16#0D#),
      2572 => to_slv(opcode_type, 16#0D#),
      2573 => to_slv(opcode_type, 16#06#),
      2574 => to_slv(opcode_type, 16#10#),
      2575 => to_slv(opcode_type, 16#0C#),
      2576 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#03#),
      2593 => to_slv(opcode_type, 16#08#),
      2594 => to_slv(opcode_type, 16#07#),
      2595 => to_slv(opcode_type, 16#09#),
      2596 => to_slv(opcode_type, 16#11#),
      2597 => to_slv(opcode_type, 16#11#),
      2598 => to_slv(opcode_type, 16#09#),
      2599 => to_slv(opcode_type, 16#0A#),
      2600 => to_slv(opcode_type, 16#0F#),
      2601 => to_slv(opcode_type, 16#08#),
      2602 => to_slv(opcode_type, 16#08#),
      2603 => to_slv(opcode_type, 16#0A#),
      2604 => to_slv(opcode_type, 16#0A#),
      2605 => to_slv(opcode_type, 16#07#),
      2606 => to_slv(opcode_type, 16#10#),
      2607 => to_slv(opcode_type, 16#0D#),
      2608 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#09#),
      2625 => to_slv(opcode_type, 16#06#),
      2626 => to_slv(opcode_type, 16#06#),
      2627 => to_slv(opcode_type, 16#09#),
      2628 => to_slv(opcode_type, 16#0C#),
      2629 => to_slv(opcode_type, 16#0D#),
      2630 => to_slv(opcode_type, 16#05#),
      2631 => to_slv(opcode_type, 16#0B#),
      2632 => to_slv(opcode_type, 16#07#),
      2633 => to_slv(opcode_type, 16#01#),
      2634 => to_slv(opcode_type, 16#68#),
      2635 => to_slv(opcode_type, 16#08#),
      2636 => to_slv(opcode_type, 16#0C#),
      2637 => to_slv(opcode_type, 16#0D#),
      2638 => to_slv(opcode_type, 16#05#),
      2639 => to_slv(opcode_type, 16#11#),
      2640 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#09#),
      2657 => to_slv(opcode_type, 16#02#),
      2658 => to_slv(opcode_type, 16#03#),
      2659 => to_slv(opcode_type, 16#02#),
      2660 => to_slv(opcode_type, 16#0C#),
      2661 => to_slv(opcode_type, 16#06#),
      2662 => to_slv(opcode_type, 16#04#),
      2663 => to_slv(opcode_type, 16#07#),
      2664 => to_slv(opcode_type, 16#0D#),
      2665 => to_slv(opcode_type, 16#0A#),
      2666 => to_slv(opcode_type, 16#08#),
      2667 => to_slv(opcode_type, 16#08#),
      2668 => to_slv(opcode_type, 16#10#),
      2669 => to_slv(opcode_type, 16#10#),
      2670 => to_slv(opcode_type, 16#03#),
      2671 => to_slv(opcode_type, 16#0E#),
      2672 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#04#),
      2689 => to_slv(opcode_type, 16#09#),
      2690 => to_slv(opcode_type, 16#07#),
      2691 => to_slv(opcode_type, 16#08#),
      2692 => to_slv(opcode_type, 16#0B#),
      2693 => to_slv(opcode_type, 16#0A#),
      2694 => to_slv(opcode_type, 16#09#),
      2695 => to_slv(opcode_type, 16#0E#),
      2696 => to_slv(opcode_type, 16#F8#),
      2697 => to_slv(opcode_type, 16#06#),
      2698 => to_slv(opcode_type, 16#06#),
      2699 => to_slv(opcode_type, 16#0E#),
      2700 => to_slv(opcode_type, 16#0B#),
      2701 => to_slv(opcode_type, 16#08#),
      2702 => to_slv(opcode_type, 16#0F#),
      2703 => to_slv(opcode_type, 16#0C#),
      2704 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#03#),
      2721 => to_slv(opcode_type, 16#08#),
      2722 => to_slv(opcode_type, 16#08#),
      2723 => to_slv(opcode_type, 16#08#),
      2724 => to_slv(opcode_type, 16#0D#),
      2725 => to_slv(opcode_type, 16#0B#),
      2726 => to_slv(opcode_type, 16#06#),
      2727 => to_slv(opcode_type, 16#B9#),
      2728 => to_slv(opcode_type, 16#0F#),
      2729 => to_slv(opcode_type, 16#08#),
      2730 => to_slv(opcode_type, 16#06#),
      2731 => to_slv(opcode_type, 16#0B#),
      2732 => to_slv(opcode_type, 16#0D#),
      2733 => to_slv(opcode_type, 16#08#),
      2734 => to_slv(opcode_type, 16#0D#),
      2735 => to_slv(opcode_type, 16#11#),
      2736 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#09#),
      2753 => to_slv(opcode_type, 16#07#),
      2754 => to_slv(opcode_type, 16#08#),
      2755 => to_slv(opcode_type, 16#08#),
      2756 => to_slv(opcode_type, 16#0B#),
      2757 => to_slv(opcode_type, 16#0B#),
      2758 => to_slv(opcode_type, 16#07#),
      2759 => to_slv(opcode_type, 16#0D#),
      2760 => to_slv(opcode_type, 16#11#),
      2761 => to_slv(opcode_type, 16#04#),
      2762 => to_slv(opcode_type, 16#08#),
      2763 => to_slv(opcode_type, 16#10#),
      2764 => to_slv(opcode_type, 16#0C#),
      2765 => to_slv(opcode_type, 16#07#),
      2766 => to_slv(opcode_type, 16#0E#),
      2767 => to_slv(opcode_type, 16#10#),
      2768 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#08#),
      2785 => to_slv(opcode_type, 16#05#),
      2786 => to_slv(opcode_type, 16#01#),
      2787 => to_slv(opcode_type, 16#07#),
      2788 => to_slv(opcode_type, 16#0F#),
      2789 => to_slv(opcode_type, 16#0F#),
      2790 => to_slv(opcode_type, 16#09#),
      2791 => to_slv(opcode_type, 16#03#),
      2792 => to_slv(opcode_type, 16#09#),
      2793 => to_slv(opcode_type, 16#0B#),
      2794 => to_slv(opcode_type, 16#0C#),
      2795 => to_slv(opcode_type, 16#06#),
      2796 => to_slv(opcode_type, 16#07#),
      2797 => to_slv(opcode_type, 16#1C#),
      2798 => to_slv(opcode_type, 16#49#),
      2799 => to_slv(opcode_type, 16#B1#),
      2800 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#04#),
      2817 => to_slv(opcode_type, 16#09#),
      2818 => to_slv(opcode_type, 16#09#),
      2819 => to_slv(opcode_type, 16#09#),
      2820 => to_slv(opcode_type, 16#0E#),
      2821 => to_slv(opcode_type, 16#0E#),
      2822 => to_slv(opcode_type, 16#06#),
      2823 => to_slv(opcode_type, 16#0F#),
      2824 => to_slv(opcode_type, 16#11#),
      2825 => to_slv(opcode_type, 16#07#),
      2826 => to_slv(opcode_type, 16#06#),
      2827 => to_slv(opcode_type, 16#0D#),
      2828 => to_slv(opcode_type, 16#0D#),
      2829 => to_slv(opcode_type, 16#09#),
      2830 => to_slv(opcode_type, 16#0E#),
      2831 => to_slv(opcode_type, 16#0F#),
      2832 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#09#),
      2849 => to_slv(opcode_type, 16#01#),
      2850 => to_slv(opcode_type, 16#06#),
      2851 => to_slv(opcode_type, 16#04#),
      2852 => to_slv(opcode_type, 16#11#),
      2853 => to_slv(opcode_type, 16#06#),
      2854 => to_slv(opcode_type, 16#0A#),
      2855 => to_slv(opcode_type, 16#0E#),
      2856 => to_slv(opcode_type, 16#08#),
      2857 => to_slv(opcode_type, 16#04#),
      2858 => to_slv(opcode_type, 16#02#),
      2859 => to_slv(opcode_type, 16#0D#),
      2860 => to_slv(opcode_type, 16#08#),
      2861 => to_slv(opcode_type, 16#01#),
      2862 => to_slv(opcode_type, 16#5A#),
      2863 => to_slv(opcode_type, 16#0C#),
      2864 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#01#),
      2881 => to_slv(opcode_type, 16#06#),
      2882 => to_slv(opcode_type, 16#06#),
      2883 => to_slv(opcode_type, 16#06#),
      2884 => to_slv(opcode_type, 16#0C#),
      2885 => to_slv(opcode_type, 16#0F#),
      2886 => to_slv(opcode_type, 16#07#),
      2887 => to_slv(opcode_type, 16#0E#),
      2888 => to_slv(opcode_type, 16#10#),
      2889 => to_slv(opcode_type, 16#09#),
      2890 => to_slv(opcode_type, 16#09#),
      2891 => to_slv(opcode_type, 16#87#),
      2892 => to_slv(opcode_type, 16#10#),
      2893 => to_slv(opcode_type, 16#07#),
      2894 => to_slv(opcode_type, 16#10#),
      2895 => to_slv(opcode_type, 16#11#),
      2896 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#09#),
      2913 => to_slv(opcode_type, 16#03#),
      2914 => to_slv(opcode_type, 16#05#),
      2915 => to_slv(opcode_type, 16#05#),
      2916 => to_slv(opcode_type, 16#0B#),
      2917 => to_slv(opcode_type, 16#09#),
      2918 => to_slv(opcode_type, 16#08#),
      2919 => to_slv(opcode_type, 16#08#),
      2920 => to_slv(opcode_type, 16#0A#),
      2921 => to_slv(opcode_type, 16#0B#),
      2922 => to_slv(opcode_type, 16#04#),
      2923 => to_slv(opcode_type, 16#10#),
      2924 => to_slv(opcode_type, 16#01#),
      2925 => to_slv(opcode_type, 16#08#),
      2926 => to_slv(opcode_type, 16#0D#),
      2927 => to_slv(opcode_type, 16#0D#),
      2928 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#09#),
      2945 => to_slv(opcode_type, 16#01#),
      2946 => to_slv(opcode_type, 16#06#),
      2947 => to_slv(opcode_type, 16#04#),
      2948 => to_slv(opcode_type, 16#7E#),
      2949 => to_slv(opcode_type, 16#01#),
      2950 => to_slv(opcode_type, 16#0F#),
      2951 => to_slv(opcode_type, 16#09#),
      2952 => to_slv(opcode_type, 16#03#),
      2953 => to_slv(opcode_type, 16#08#),
      2954 => to_slv(opcode_type, 16#0C#),
      2955 => to_slv(opcode_type, 16#0C#),
      2956 => to_slv(opcode_type, 16#02#),
      2957 => to_slv(opcode_type, 16#09#),
      2958 => to_slv(opcode_type, 16#0A#),
      2959 => to_slv(opcode_type, 16#0C#),
      2960 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#04#),
      2977 => to_slv(opcode_type, 16#07#),
      2978 => to_slv(opcode_type, 16#09#),
      2979 => to_slv(opcode_type, 16#08#),
      2980 => to_slv(opcode_type, 16#0D#),
      2981 => to_slv(opcode_type, 16#B9#),
      2982 => to_slv(opcode_type, 16#08#),
      2983 => to_slv(opcode_type, 16#11#),
      2984 => to_slv(opcode_type, 16#0A#),
      2985 => to_slv(opcode_type, 16#06#),
      2986 => to_slv(opcode_type, 16#07#),
      2987 => to_slv(opcode_type, 16#0F#),
      2988 => to_slv(opcode_type, 16#10#),
      2989 => to_slv(opcode_type, 16#06#),
      2990 => to_slv(opcode_type, 16#57#),
      2991 => to_slv(opcode_type, 16#0D#),
      2992 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#04#),
      3009 => to_slv(opcode_type, 16#08#),
      3010 => to_slv(opcode_type, 16#07#),
      3011 => to_slv(opcode_type, 16#07#),
      3012 => to_slv(opcode_type, 16#11#),
      3013 => to_slv(opcode_type, 16#0A#),
      3014 => to_slv(opcode_type, 16#08#),
      3015 => to_slv(opcode_type, 16#0F#),
      3016 => to_slv(opcode_type, 16#0A#),
      3017 => to_slv(opcode_type, 16#08#),
      3018 => to_slv(opcode_type, 16#07#),
      3019 => to_slv(opcode_type, 16#0E#),
      3020 => to_slv(opcode_type, 16#0F#),
      3021 => to_slv(opcode_type, 16#06#),
      3022 => to_slv(opcode_type, 16#11#),
      3023 => to_slv(opcode_type, 16#0E#),
      3024 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#03#),
      3041 => to_slv(opcode_type, 16#06#),
      3042 => to_slv(opcode_type, 16#09#),
      3043 => to_slv(opcode_type, 16#06#),
      3044 => to_slv(opcode_type, 16#0E#),
      3045 => to_slv(opcode_type, 16#0F#),
      3046 => to_slv(opcode_type, 16#08#),
      3047 => to_slv(opcode_type, 16#0D#),
      3048 => to_slv(opcode_type, 16#10#),
      3049 => to_slv(opcode_type, 16#08#),
      3050 => to_slv(opcode_type, 16#07#),
      3051 => to_slv(opcode_type, 16#0B#),
      3052 => to_slv(opcode_type, 16#0B#),
      3053 => to_slv(opcode_type, 16#08#),
      3054 => to_slv(opcode_type, 16#0F#),
      3055 => to_slv(opcode_type, 16#0F#),
      3056 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#05#),
      3073 => to_slv(opcode_type, 16#09#),
      3074 => to_slv(opcode_type, 16#08#),
      3075 => to_slv(opcode_type, 16#08#),
      3076 => to_slv(opcode_type, 16#0C#),
      3077 => to_slv(opcode_type, 16#0A#),
      3078 => to_slv(opcode_type, 16#09#),
      3079 => to_slv(opcode_type, 16#0B#),
      3080 => to_slv(opcode_type, 16#0D#),
      3081 => to_slv(opcode_type, 16#09#),
      3082 => to_slv(opcode_type, 16#07#),
      3083 => to_slv(opcode_type, 16#0E#),
      3084 => to_slv(opcode_type, 16#0C#),
      3085 => to_slv(opcode_type, 16#07#),
      3086 => to_slv(opcode_type, 16#11#),
      3087 => to_slv(opcode_type, 16#10#),
      3088 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#06#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#02#),
      3107 => to_slv(opcode_type, 16#03#),
      3108 => to_slv(opcode_type, 16#0E#),
      3109 => to_slv(opcode_type, 16#02#),
      3110 => to_slv(opcode_type, 16#09#),
      3111 => to_slv(opcode_type, 16#0B#),
      3112 => to_slv(opcode_type, 16#0E#),
      3113 => to_slv(opcode_type, 16#02#),
      3114 => to_slv(opcode_type, 16#07#),
      3115 => to_slv(opcode_type, 16#07#),
      3116 => to_slv(opcode_type, 16#0A#),
      3117 => to_slv(opcode_type, 16#0D#),
      3118 => to_slv(opcode_type, 16#04#),
      3119 => to_slv(opcode_type, 16#0C#),
      3120 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#03#),
      3137 => to_slv(opcode_type, 16#08#),
      3138 => to_slv(opcode_type, 16#06#),
      3139 => to_slv(opcode_type, 16#06#),
      3140 => to_slv(opcode_type, 16#11#),
      3141 => to_slv(opcode_type, 16#0B#),
      3142 => to_slv(opcode_type, 16#07#),
      3143 => to_slv(opcode_type, 16#10#),
      3144 => to_slv(opcode_type, 16#0F#),
      3145 => to_slv(opcode_type, 16#08#),
      3146 => to_slv(opcode_type, 16#08#),
      3147 => to_slv(opcode_type, 16#0B#),
      3148 => to_slv(opcode_type, 16#0D#),
      3149 => to_slv(opcode_type, 16#06#),
      3150 => to_slv(opcode_type, 16#0A#),
      3151 => to_slv(opcode_type, 16#10#),
      3152 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#03#),
      3169 => to_slv(opcode_type, 16#09#),
      3170 => to_slv(opcode_type, 16#09#),
      3171 => to_slv(opcode_type, 16#07#),
      3172 => to_slv(opcode_type, 16#0F#),
      3173 => to_slv(opcode_type, 16#0C#),
      3174 => to_slv(opcode_type, 16#07#),
      3175 => to_slv(opcode_type, 16#0B#),
      3176 => to_slv(opcode_type, 16#0C#),
      3177 => to_slv(opcode_type, 16#09#),
      3178 => to_slv(opcode_type, 16#07#),
      3179 => to_slv(opcode_type, 16#0E#),
      3180 => to_slv(opcode_type, 16#85#),
      3181 => to_slv(opcode_type, 16#06#),
      3182 => to_slv(opcode_type, 16#0F#),
      3183 => to_slv(opcode_type, 16#10#),
      3184 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#06#),
      3201 => to_slv(opcode_type, 16#01#),
      3202 => to_slv(opcode_type, 16#06#),
      3203 => to_slv(opcode_type, 16#02#),
      3204 => to_slv(opcode_type, 16#0D#),
      3205 => to_slv(opcode_type, 16#05#),
      3206 => to_slv(opcode_type, 16#0F#),
      3207 => to_slv(opcode_type, 16#08#),
      3208 => to_slv(opcode_type, 16#09#),
      3209 => to_slv(opcode_type, 16#09#),
      3210 => to_slv(opcode_type, 16#11#),
      3211 => to_slv(opcode_type, 16#0B#),
      3212 => to_slv(opcode_type, 16#05#),
      3213 => to_slv(opcode_type, 16#0D#),
      3214 => to_slv(opcode_type, 16#04#),
      3215 => to_slv(opcode_type, 16#0A#),
      3216 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#03#),
      3233 => to_slv(opcode_type, 16#08#),
      3234 => to_slv(opcode_type, 16#08#),
      3235 => to_slv(opcode_type, 16#09#),
      3236 => to_slv(opcode_type, 16#0B#),
      3237 => to_slv(opcode_type, 16#0F#),
      3238 => to_slv(opcode_type, 16#08#),
      3239 => to_slv(opcode_type, 16#10#),
      3240 => to_slv(opcode_type, 16#0F#),
      3241 => to_slv(opcode_type, 16#06#),
      3242 => to_slv(opcode_type, 16#08#),
      3243 => to_slv(opcode_type, 16#10#),
      3244 => to_slv(opcode_type, 16#10#),
      3245 => to_slv(opcode_type, 16#09#),
      3246 => to_slv(opcode_type, 16#11#),
      3247 => to_slv(opcode_type, 16#0D#),
      3248 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#09#),
      3265 => to_slv(opcode_type, 16#07#),
      3266 => to_slv(opcode_type, 16#02#),
      3267 => to_slv(opcode_type, 16#04#),
      3268 => to_slv(opcode_type, 16#0D#),
      3269 => to_slv(opcode_type, 16#09#),
      3270 => to_slv(opcode_type, 16#03#),
      3271 => to_slv(opcode_type, 16#11#),
      3272 => to_slv(opcode_type, 16#06#),
      3273 => to_slv(opcode_type, 16#0C#),
      3274 => to_slv(opcode_type, 16#0D#),
      3275 => to_slv(opcode_type, 16#09#),
      3276 => to_slv(opcode_type, 16#09#),
      3277 => to_slv(opcode_type, 16#0E#),
      3278 => to_slv(opcode_type, 16#0D#),
      3279 => to_slv(opcode_type, 16#10#),
      3280 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#08#),
      3297 => to_slv(opcode_type, 16#01#),
      3298 => to_slv(opcode_type, 16#04#),
      3299 => to_slv(opcode_type, 16#07#),
      3300 => to_slv(opcode_type, 16#0C#),
      3301 => to_slv(opcode_type, 16#0B#),
      3302 => to_slv(opcode_type, 16#09#),
      3303 => to_slv(opcode_type, 16#05#),
      3304 => to_slv(opcode_type, 16#03#),
      3305 => to_slv(opcode_type, 16#0E#),
      3306 => to_slv(opcode_type, 16#09#),
      3307 => to_slv(opcode_type, 16#02#),
      3308 => to_slv(opcode_type, 16#51#),
      3309 => to_slv(opcode_type, 16#09#),
      3310 => to_slv(opcode_type, 16#0F#),
      3311 => to_slv(opcode_type, 16#10#),
      3312 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#02#),
      3329 => to_slv(opcode_type, 16#08#),
      3330 => to_slv(opcode_type, 16#07#),
      3331 => to_slv(opcode_type, 16#09#),
      3332 => to_slv(opcode_type, 16#81#),
      3333 => to_slv(opcode_type, 16#0F#),
      3334 => to_slv(opcode_type, 16#06#),
      3335 => to_slv(opcode_type, 16#10#),
      3336 => to_slv(opcode_type, 16#0A#),
      3337 => to_slv(opcode_type, 16#06#),
      3338 => to_slv(opcode_type, 16#06#),
      3339 => to_slv(opcode_type, 16#0B#),
      3340 => to_slv(opcode_type, 16#0A#),
      3341 => to_slv(opcode_type, 16#09#),
      3342 => to_slv(opcode_type, 16#0E#),
      3343 => to_slv(opcode_type, 16#0A#),
      3344 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#02#),
      3361 => to_slv(opcode_type, 16#07#),
      3362 => to_slv(opcode_type, 16#07#),
      3363 => to_slv(opcode_type, 16#07#),
      3364 => to_slv(opcode_type, 16#0D#),
      3365 => to_slv(opcode_type, 16#0F#),
      3366 => to_slv(opcode_type, 16#07#),
      3367 => to_slv(opcode_type, 16#0E#),
      3368 => to_slv(opcode_type, 16#0C#),
      3369 => to_slv(opcode_type, 16#07#),
      3370 => to_slv(opcode_type, 16#06#),
      3371 => to_slv(opcode_type, 16#0E#),
      3372 => to_slv(opcode_type, 16#0A#),
      3373 => to_slv(opcode_type, 16#08#),
      3374 => to_slv(opcode_type, 16#10#),
      3375 => to_slv(opcode_type, 16#0F#),
      3376 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#08#),
      3393 => to_slv(opcode_type, 16#04#),
      3394 => to_slv(opcode_type, 16#07#),
      3395 => to_slv(opcode_type, 16#01#),
      3396 => to_slv(opcode_type, 16#57#),
      3397 => to_slv(opcode_type, 16#04#),
      3398 => to_slv(opcode_type, 16#11#),
      3399 => to_slv(opcode_type, 16#08#),
      3400 => to_slv(opcode_type, 16#03#),
      3401 => to_slv(opcode_type, 16#06#),
      3402 => to_slv(opcode_type, 16#0B#),
      3403 => to_slv(opcode_type, 16#0F#),
      3404 => to_slv(opcode_type, 16#02#),
      3405 => to_slv(opcode_type, 16#08#),
      3406 => to_slv(opcode_type, 16#0B#),
      3407 => to_slv(opcode_type, 16#0B#),
      3408 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#03#),
      3426 => to_slv(opcode_type, 16#02#),
      3427 => to_slv(opcode_type, 16#04#),
      3428 => to_slv(opcode_type, 16#0C#),
      3429 => to_slv(opcode_type, 16#09#),
      3430 => to_slv(opcode_type, 16#09#),
      3431 => to_slv(opcode_type, 16#06#),
      3432 => to_slv(opcode_type, 16#11#),
      3433 => to_slv(opcode_type, 16#11#),
      3434 => to_slv(opcode_type, 16#07#),
      3435 => to_slv(opcode_type, 16#10#),
      3436 => to_slv(opcode_type, 16#11#),
      3437 => to_slv(opcode_type, 16#08#),
      3438 => to_slv(opcode_type, 16#10#),
      3439 => to_slv(opcode_type, 16#0F#),
      3440 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#05#),
      3457 => to_slv(opcode_type, 16#06#),
      3458 => to_slv(opcode_type, 16#08#),
      3459 => to_slv(opcode_type, 16#09#),
      3460 => to_slv(opcode_type, 16#0F#),
      3461 => to_slv(opcode_type, 16#11#),
      3462 => to_slv(opcode_type, 16#06#),
      3463 => to_slv(opcode_type, 16#0E#),
      3464 => to_slv(opcode_type, 16#0E#),
      3465 => to_slv(opcode_type, 16#07#),
      3466 => to_slv(opcode_type, 16#06#),
      3467 => to_slv(opcode_type, 16#0A#),
      3468 => to_slv(opcode_type, 16#0D#),
      3469 => to_slv(opcode_type, 16#09#),
      3470 => to_slv(opcode_type, 16#11#),
      3471 => to_slv(opcode_type, 16#0C#),
      3472 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#09#),
      3489 => to_slv(opcode_type, 16#07#),
      3490 => to_slv(opcode_type, 16#03#),
      3491 => to_slv(opcode_type, 16#07#),
      3492 => to_slv(opcode_type, 16#10#),
      3493 => to_slv(opcode_type, 16#0D#),
      3494 => to_slv(opcode_type, 16#08#),
      3495 => to_slv(opcode_type, 16#05#),
      3496 => to_slv(opcode_type, 16#10#),
      3497 => to_slv(opcode_type, 16#07#),
      3498 => to_slv(opcode_type, 16#0D#),
      3499 => to_slv(opcode_type, 16#0B#),
      3500 => to_slv(opcode_type, 16#01#),
      3501 => to_slv(opcode_type, 16#04#),
      3502 => to_slv(opcode_type, 16#01#),
      3503 => to_slv(opcode_type, 16#0D#),
      3504 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#08#),
      3521 => to_slv(opcode_type, 16#06#),
      3522 => to_slv(opcode_type, 16#03#),
      3523 => to_slv(opcode_type, 16#05#),
      3524 => to_slv(opcode_type, 16#0A#),
      3525 => to_slv(opcode_type, 16#09#),
      3526 => to_slv(opcode_type, 16#09#),
      3527 => to_slv(opcode_type, 16#0E#),
      3528 => to_slv(opcode_type, 16#11#),
      3529 => to_slv(opcode_type, 16#04#),
      3530 => to_slv(opcode_type, 16#11#),
      3531 => to_slv(opcode_type, 16#09#),
      3532 => to_slv(opcode_type, 16#03#),
      3533 => to_slv(opcode_type, 16#04#),
      3534 => to_slv(opcode_type, 16#11#),
      3535 => to_slv(opcode_type, 16#10#),
      3536 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#07#),
      3553 => to_slv(opcode_type, 16#01#),
      3554 => to_slv(opcode_type, 16#09#),
      3555 => to_slv(opcode_type, 16#01#),
      3556 => to_slv(opcode_type, 16#0A#),
      3557 => to_slv(opcode_type, 16#08#),
      3558 => to_slv(opcode_type, 16#10#),
      3559 => to_slv(opcode_type, 16#0F#),
      3560 => to_slv(opcode_type, 16#07#),
      3561 => to_slv(opcode_type, 16#05#),
      3562 => to_slv(opcode_type, 16#02#),
      3563 => to_slv(opcode_type, 16#0D#),
      3564 => to_slv(opcode_type, 16#03#),
      3565 => to_slv(opcode_type, 16#09#),
      3566 => to_slv(opcode_type, 16#0F#),
      3567 => to_slv(opcode_type, 16#0E#),
      3568 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#03#),
      3585 => to_slv(opcode_type, 16#06#),
      3586 => to_slv(opcode_type, 16#07#),
      3587 => to_slv(opcode_type, 16#08#),
      3588 => to_slv(opcode_type, 16#11#),
      3589 => to_slv(opcode_type, 16#0A#),
      3590 => to_slv(opcode_type, 16#07#),
      3591 => to_slv(opcode_type, 16#11#),
      3592 => to_slv(opcode_type, 16#0D#),
      3593 => to_slv(opcode_type, 16#06#),
      3594 => to_slv(opcode_type, 16#07#),
      3595 => to_slv(opcode_type, 16#11#),
      3596 => to_slv(opcode_type, 16#0F#),
      3597 => to_slv(opcode_type, 16#06#),
      3598 => to_slv(opcode_type, 16#0E#),
      3599 => to_slv(opcode_type, 16#11#),
      3600 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#01#),
      3617 => to_slv(opcode_type, 16#09#),
      3618 => to_slv(opcode_type, 16#09#),
      3619 => to_slv(opcode_type, 16#06#),
      3620 => to_slv(opcode_type, 16#10#),
      3621 => to_slv(opcode_type, 16#0A#),
      3622 => to_slv(opcode_type, 16#07#),
      3623 => to_slv(opcode_type, 16#0E#),
      3624 => to_slv(opcode_type, 16#0D#),
      3625 => to_slv(opcode_type, 16#08#),
      3626 => to_slv(opcode_type, 16#07#),
      3627 => to_slv(opcode_type, 16#0F#),
      3628 => to_slv(opcode_type, 16#33#),
      3629 => to_slv(opcode_type, 16#08#),
      3630 => to_slv(opcode_type, 16#11#),
      3631 => to_slv(opcode_type, 16#0C#),
      3632 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#07#),
      3649 => to_slv(opcode_type, 16#09#),
      3650 => to_slv(opcode_type, 16#03#),
      3651 => to_slv(opcode_type, 16#02#),
      3652 => to_slv(opcode_type, 16#0B#),
      3653 => to_slv(opcode_type, 16#02#),
      3654 => to_slv(opcode_type, 16#09#),
      3655 => to_slv(opcode_type, 16#0A#),
      3656 => to_slv(opcode_type, 16#0B#),
      3657 => to_slv(opcode_type, 16#08#),
      3658 => to_slv(opcode_type, 16#06#),
      3659 => to_slv(opcode_type, 16#05#),
      3660 => to_slv(opcode_type, 16#10#),
      3661 => to_slv(opcode_type, 16#04#),
      3662 => to_slv(opcode_type, 16#0D#),
      3663 => to_slv(opcode_type, 16#0B#),
      3664 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#01#),
      3681 => to_slv(opcode_type, 16#09#),
      3682 => to_slv(opcode_type, 16#06#),
      3683 => to_slv(opcode_type, 16#08#),
      3684 => to_slv(opcode_type, 16#0C#),
      3685 => to_slv(opcode_type, 16#10#),
      3686 => to_slv(opcode_type, 16#09#),
      3687 => to_slv(opcode_type, 16#0F#),
      3688 => to_slv(opcode_type, 16#0F#),
      3689 => to_slv(opcode_type, 16#09#),
      3690 => to_slv(opcode_type, 16#07#),
      3691 => to_slv(opcode_type, 16#0C#),
      3692 => to_slv(opcode_type, 16#0D#),
      3693 => to_slv(opcode_type, 16#07#),
      3694 => to_slv(opcode_type, 16#0E#),
      3695 => to_slv(opcode_type, 16#0E#),
      3696 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#07#),
      3713 => to_slv(opcode_type, 16#05#),
      3714 => to_slv(opcode_type, 16#03#),
      3715 => to_slv(opcode_type, 16#02#),
      3716 => to_slv(opcode_type, 16#0F#),
      3717 => to_slv(opcode_type, 16#09#),
      3718 => to_slv(opcode_type, 16#04#),
      3719 => to_slv(opcode_type, 16#08#),
      3720 => to_slv(opcode_type, 16#9D#),
      3721 => to_slv(opcode_type, 16#0D#),
      3722 => to_slv(opcode_type, 16#06#),
      3723 => to_slv(opcode_type, 16#08#),
      3724 => to_slv(opcode_type, 16#0A#),
      3725 => to_slv(opcode_type, 16#0C#),
      3726 => to_slv(opcode_type, 16#03#),
      3727 => to_slv(opcode_type, 16#11#),
      3728 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#07#),
      3745 => to_slv(opcode_type, 16#01#),
      3746 => to_slv(opcode_type, 16#05#),
      3747 => to_slv(opcode_type, 16#03#),
      3748 => to_slv(opcode_type, 16#0D#),
      3749 => to_slv(opcode_type, 16#08#),
      3750 => to_slv(opcode_type, 16#06#),
      3751 => to_slv(opcode_type, 16#06#),
      3752 => to_slv(opcode_type, 16#0B#),
      3753 => to_slv(opcode_type, 16#0A#),
      3754 => to_slv(opcode_type, 16#05#),
      3755 => to_slv(opcode_type, 16#E7#),
      3756 => to_slv(opcode_type, 16#07#),
      3757 => to_slv(opcode_type, 16#01#),
      3758 => to_slv(opcode_type, 16#0C#),
      3759 => to_slv(opcode_type, 16#0C#),
      3760 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#07#),
      3777 => to_slv(opcode_type, 16#06#),
      3778 => to_slv(opcode_type, 16#02#),
      3779 => to_slv(opcode_type, 16#05#),
      3780 => to_slv(opcode_type, 16#0A#),
      3781 => to_slv(opcode_type, 16#01#),
      3782 => to_slv(opcode_type, 16#08#),
      3783 => to_slv(opcode_type, 16#0E#),
      3784 => to_slv(opcode_type, 16#0C#),
      3785 => to_slv(opcode_type, 16#09#),
      3786 => to_slv(opcode_type, 16#06#),
      3787 => to_slv(opcode_type, 16#04#),
      3788 => to_slv(opcode_type, 16#0C#),
      3789 => to_slv(opcode_type, 16#05#),
      3790 => to_slv(opcode_type, 16#10#),
      3791 => to_slv(opcode_type, 16#0A#),
      3792 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#04#),
      3809 => to_slv(opcode_type, 16#07#),
      3810 => to_slv(opcode_type, 16#06#),
      3811 => to_slv(opcode_type, 16#08#),
      3812 => to_slv(opcode_type, 16#0B#),
      3813 => to_slv(opcode_type, 16#0A#),
      3814 => to_slv(opcode_type, 16#06#),
      3815 => to_slv(opcode_type, 16#0E#),
      3816 => to_slv(opcode_type, 16#0F#),
      3817 => to_slv(opcode_type, 16#07#),
      3818 => to_slv(opcode_type, 16#07#),
      3819 => to_slv(opcode_type, 16#11#),
      3820 => to_slv(opcode_type, 16#0B#),
      3821 => to_slv(opcode_type, 16#06#),
      3822 => to_slv(opcode_type, 16#0F#),
      3823 => to_slv(opcode_type, 16#11#),
      3824 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#08#),
      3841 => to_slv(opcode_type, 16#02#),
      3842 => to_slv(opcode_type, 16#03#),
      3843 => to_slv(opcode_type, 16#04#),
      3844 => to_slv(opcode_type, 16#10#),
      3845 => to_slv(opcode_type, 16#07#),
      3846 => to_slv(opcode_type, 16#07#),
      3847 => to_slv(opcode_type, 16#09#),
      3848 => to_slv(opcode_type, 16#5B#),
      3849 => to_slv(opcode_type, 16#0C#),
      3850 => to_slv(opcode_type, 16#06#),
      3851 => to_slv(opcode_type, 16#0C#),
      3852 => to_slv(opcode_type, 16#11#),
      3853 => to_slv(opcode_type, 16#05#),
      3854 => to_slv(opcode_type, 16#01#),
      3855 => to_slv(opcode_type, 16#0C#),
      3856 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#06#),
      3873 => to_slv(opcode_type, 16#08#),
      3874 => to_slv(opcode_type, 16#06#),
      3875 => to_slv(opcode_type, 16#07#),
      3876 => to_slv(opcode_type, 16#0D#),
      3877 => to_slv(opcode_type, 16#0E#),
      3878 => to_slv(opcode_type, 16#02#),
      3879 => to_slv(opcode_type, 16#34#),
      3880 => to_slv(opcode_type, 16#02#),
      3881 => to_slv(opcode_type, 16#04#),
      3882 => to_slv(opcode_type, 16#10#),
      3883 => to_slv(opcode_type, 16#01#),
      3884 => to_slv(opcode_type, 16#08#),
      3885 => to_slv(opcode_type, 16#05#),
      3886 => to_slv(opcode_type, 16#9D#),
      3887 => to_slv(opcode_type, 16#0D#),
      3888 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#08#),
      3905 => to_slv(opcode_type, 16#02#),
      3906 => to_slv(opcode_type, 16#05#),
      3907 => to_slv(opcode_type, 16#01#),
      3908 => to_slv(opcode_type, 16#10#),
      3909 => to_slv(opcode_type, 16#08#),
      3910 => to_slv(opcode_type, 16#08#),
      3911 => to_slv(opcode_type, 16#04#),
      3912 => to_slv(opcode_type, 16#0C#),
      3913 => to_slv(opcode_type, 16#07#),
      3914 => to_slv(opcode_type, 16#0A#),
      3915 => to_slv(opcode_type, 16#9E#),
      3916 => to_slv(opcode_type, 16#02#),
      3917 => to_slv(opcode_type, 16#06#),
      3918 => to_slv(opcode_type, 16#0E#),
      3919 => to_slv(opcode_type, 16#0E#),
      3920 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#03#),
      3937 => to_slv(opcode_type, 16#08#),
      3938 => to_slv(opcode_type, 16#07#),
      3939 => to_slv(opcode_type, 16#09#),
      3940 => to_slv(opcode_type, 16#0C#),
      3941 => to_slv(opcode_type, 16#0A#),
      3942 => to_slv(opcode_type, 16#08#),
      3943 => to_slv(opcode_type, 16#0C#),
      3944 => to_slv(opcode_type, 16#0F#),
      3945 => to_slv(opcode_type, 16#09#),
      3946 => to_slv(opcode_type, 16#09#),
      3947 => to_slv(opcode_type, 16#0D#),
      3948 => to_slv(opcode_type, 16#0F#),
      3949 => to_slv(opcode_type, 16#06#),
      3950 => to_slv(opcode_type, 16#0D#),
      3951 => to_slv(opcode_type, 16#0E#),
      3952 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#08#),
      3969 => to_slv(opcode_type, 16#01#),
      3970 => to_slv(opcode_type, 16#02#),
      3971 => to_slv(opcode_type, 16#03#),
      3972 => to_slv(opcode_type, 16#0D#),
      3973 => to_slv(opcode_type, 16#09#),
      3974 => to_slv(opcode_type, 16#06#),
      3975 => to_slv(opcode_type, 16#09#),
      3976 => to_slv(opcode_type, 16#0A#),
      3977 => to_slv(opcode_type, 16#0C#),
      3978 => to_slv(opcode_type, 16#02#),
      3979 => to_slv(opcode_type, 16#0B#),
      3980 => to_slv(opcode_type, 16#01#),
      3981 => to_slv(opcode_type, 16#07#),
      3982 => to_slv(opcode_type, 16#0B#),
      3983 => to_slv(opcode_type, 16#0E#),
      3984 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#05#),
      4001 => to_slv(opcode_type, 16#08#),
      4002 => to_slv(opcode_type, 16#07#),
      4003 => to_slv(opcode_type, 16#06#),
      4004 => to_slv(opcode_type, 16#10#),
      4005 => to_slv(opcode_type, 16#0A#),
      4006 => to_slv(opcode_type, 16#08#),
      4007 => to_slv(opcode_type, 16#0F#),
      4008 => to_slv(opcode_type, 16#11#),
      4009 => to_slv(opcode_type, 16#06#),
      4010 => to_slv(opcode_type, 16#07#),
      4011 => to_slv(opcode_type, 16#AD#),
      4012 => to_slv(opcode_type, 16#0B#),
      4013 => to_slv(opcode_type, 16#07#),
      4014 => to_slv(opcode_type, 16#0E#),
      4015 => to_slv(opcode_type, 16#10#),
      4016 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#05#),
      4033 => to_slv(opcode_type, 16#07#),
      4034 => to_slv(opcode_type, 16#09#),
      4035 => to_slv(opcode_type, 16#06#),
      4036 => to_slv(opcode_type, 16#34#),
      4037 => to_slv(opcode_type, 16#10#),
      4038 => to_slv(opcode_type, 16#09#),
      4039 => to_slv(opcode_type, 16#30#),
      4040 => to_slv(opcode_type, 16#11#),
      4041 => to_slv(opcode_type, 16#06#),
      4042 => to_slv(opcode_type, 16#06#),
      4043 => to_slv(opcode_type, 16#10#),
      4044 => to_slv(opcode_type, 16#0B#),
      4045 => to_slv(opcode_type, 16#07#),
      4046 => to_slv(opcode_type, 16#0D#),
      4047 => to_slv(opcode_type, 16#10#),
      4048 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#02#),
      4066 => to_slv(opcode_type, 16#09#),
      4067 => to_slv(opcode_type, 16#06#),
      4068 => to_slv(opcode_type, 16#0A#),
      4069 => to_slv(opcode_type, 16#0F#),
      4070 => to_slv(opcode_type, 16#08#),
      4071 => to_slv(opcode_type, 16#0A#),
      4072 => to_slv(opcode_type, 16#0E#),
      4073 => to_slv(opcode_type, 16#05#),
      4074 => to_slv(opcode_type, 16#09#),
      4075 => to_slv(opcode_type, 16#05#),
      4076 => to_slv(opcode_type, 16#0B#),
      4077 => to_slv(opcode_type, 16#06#),
      4078 => to_slv(opcode_type, 16#0D#),
      4079 => to_slv(opcode_type, 16#0D#),
      4080 to 4095 => (others => '0')
  ),

    -- Bin `17`...
    16 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#06#),
      1 => to_slv(opcode_type, 16#04#),
      2 => to_slv(opcode_type, 16#02#),
      3 => to_slv(opcode_type, 16#03#),
      4 => to_slv(opcode_type, 16#0E#),
      5 => to_slv(opcode_type, 16#06#),
      6 => to_slv(opcode_type, 16#02#),
      7 => to_slv(opcode_type, 16#09#),
      8 => to_slv(opcode_type, 16#0C#),
      9 => to_slv(opcode_type, 16#0D#),
      10 => to_slv(opcode_type, 16#08#),
      11 => to_slv(opcode_type, 16#07#),
      12 => to_slv(opcode_type, 16#10#),
      13 => to_slv(opcode_type, 16#0A#),
      14 => to_slv(opcode_type, 16#09#),
      15 => to_slv(opcode_type, 16#0C#),
      16 => to_slv(opcode_type, 16#0C#),
      17 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#07#),
      33 => to_slv(opcode_type, 16#06#),
      34 => to_slv(opcode_type, 16#08#),
      35 => to_slv(opcode_type, 16#01#),
      36 => to_slv(opcode_type, 16#11#),
      37 => to_slv(opcode_type, 16#09#),
      38 => to_slv(opcode_type, 16#0C#),
      39 => to_slv(opcode_type, 16#0D#),
      40 => to_slv(opcode_type, 16#03#),
      41 => to_slv(opcode_type, 16#09#),
      42 => to_slv(opcode_type, 16#11#),
      43 => to_slv(opcode_type, 16#10#),
      44 => to_slv(opcode_type, 16#03#),
      45 => to_slv(opcode_type, 16#07#),
      46 => to_slv(opcode_type, 16#02#),
      47 => to_slv(opcode_type, 16#0F#),
      48 => to_slv(opcode_type, 16#12#),
      49 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#07#),
      65 => to_slv(opcode_type, 16#09#),
      66 => to_slv(opcode_type, 16#03#),
      67 => to_slv(opcode_type, 16#07#),
      68 => to_slv(opcode_type, 16#10#),
      69 => to_slv(opcode_type, 16#0A#),
      70 => to_slv(opcode_type, 16#08#),
      71 => to_slv(opcode_type, 16#09#),
      72 => to_slv(opcode_type, 16#0C#),
      73 => to_slv(opcode_type, 16#10#),
      74 => to_slv(opcode_type, 16#05#),
      75 => to_slv(opcode_type, 16#0C#),
      76 => to_slv(opcode_type, 16#05#),
      77 => to_slv(opcode_type, 16#04#),
      78 => to_slv(opcode_type, 16#08#),
      79 => to_slv(opcode_type, 16#0D#),
      80 => to_slv(opcode_type, 16#10#),
      81 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#06#),
      97 => to_slv(opcode_type, 16#08#),
      98 => to_slv(opcode_type, 16#07#),
      99 => to_slv(opcode_type, 16#08#),
      100 => to_slv(opcode_type, 16#0D#),
      101 => to_slv(opcode_type, 16#11#),
      102 => to_slv(opcode_type, 16#06#),
      103 => to_slv(opcode_type, 16#11#),
      104 => to_slv(opcode_type, 16#0E#),
      105 => to_slv(opcode_type, 16#05#),
      106 => to_slv(opcode_type, 16#01#),
      107 => to_slv(opcode_type, 16#0E#),
      108 => to_slv(opcode_type, 16#01#),
      109 => to_slv(opcode_type, 16#09#),
      110 => to_slv(opcode_type, 16#02#),
      111 => to_slv(opcode_type, 16#0D#),
      112 => to_slv(opcode_type, 16#87#),
      113 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#08#),
      129 => to_slv(opcode_type, 16#04#),
      130 => to_slv(opcode_type, 16#04#),
      131 => to_slv(opcode_type, 16#01#),
      132 => to_slv(opcode_type, 16#0D#),
      133 => to_slv(opcode_type, 16#09#),
      134 => to_slv(opcode_type, 16#05#),
      135 => to_slv(opcode_type, 16#09#),
      136 => to_slv(opcode_type, 16#10#),
      137 => to_slv(opcode_type, 16#10#),
      138 => to_slv(opcode_type, 16#08#),
      139 => to_slv(opcode_type, 16#06#),
      140 => to_slv(opcode_type, 16#11#),
      141 => to_slv(opcode_type, 16#0C#),
      142 => to_slv(opcode_type, 16#09#),
      143 => to_slv(opcode_type, 16#0E#),
      144 => to_slv(opcode_type, 16#0A#),
      145 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#06#),
      161 => to_slv(opcode_type, 16#03#),
      162 => to_slv(opcode_type, 16#04#),
      163 => to_slv(opcode_type, 16#02#),
      164 => to_slv(opcode_type, 16#0E#),
      165 => to_slv(opcode_type, 16#08#),
      166 => to_slv(opcode_type, 16#05#),
      167 => to_slv(opcode_type, 16#06#),
      168 => to_slv(opcode_type, 16#0B#),
      169 => to_slv(opcode_type, 16#A9#),
      170 => to_slv(opcode_type, 16#09#),
      171 => to_slv(opcode_type, 16#07#),
      172 => to_slv(opcode_type, 16#11#),
      173 => to_slv(opcode_type, 16#0A#),
      174 => to_slv(opcode_type, 16#06#),
      175 => to_slv(opcode_type, 16#0A#),
      176 => to_slv(opcode_type, 16#0D#),
      177 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#06#),
      193 => to_slv(opcode_type, 16#09#),
      194 => to_slv(opcode_type, 16#03#),
      195 => to_slv(opcode_type, 16#03#),
      196 => to_slv(opcode_type, 16#0D#),
      197 => to_slv(opcode_type, 16#03#),
      198 => to_slv(opcode_type, 16#02#),
      199 => to_slv(opcode_type, 16#0A#),
      200 => to_slv(opcode_type, 16#09#),
      201 => to_slv(opcode_type, 16#01#),
      202 => to_slv(opcode_type, 16#06#),
      203 => to_slv(opcode_type, 16#0C#),
      204 => to_slv(opcode_type, 16#0E#),
      205 => to_slv(opcode_type, 16#06#),
      206 => to_slv(opcode_type, 16#03#),
      207 => to_slv(opcode_type, 16#0B#),
      208 => to_slv(opcode_type, 16#0F#),
      209 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#07#),
      225 => to_slv(opcode_type, 16#04#),
      226 => to_slv(opcode_type, 16#06#),
      227 => to_slv(opcode_type, 16#03#),
      228 => to_slv(opcode_type, 16#11#),
      229 => to_slv(opcode_type, 16#09#),
      230 => to_slv(opcode_type, 16#0A#),
      231 => to_slv(opcode_type, 16#10#),
      232 => to_slv(opcode_type, 16#08#),
      233 => to_slv(opcode_type, 16#09#),
      234 => to_slv(opcode_type, 16#09#),
      235 => to_slv(opcode_type, 16#0A#),
      236 => to_slv(opcode_type, 16#0E#),
      237 => to_slv(opcode_type, 16#04#),
      238 => to_slv(opcode_type, 16#11#),
      239 => to_slv(opcode_type, 16#05#),
      240 => to_slv(opcode_type, 16#0A#),
      241 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#08#),
      257 => to_slv(opcode_type, 16#06#),
      258 => to_slv(opcode_type, 16#07#),
      259 => to_slv(opcode_type, 16#08#),
      260 => to_slv(opcode_type, 16#10#),
      261 => to_slv(opcode_type, 16#10#),
      262 => to_slv(opcode_type, 16#03#),
      263 => to_slv(opcode_type, 16#E6#),
      264 => to_slv(opcode_type, 16#07#),
      265 => to_slv(opcode_type, 16#02#),
      266 => to_slv(opcode_type, 16#11#),
      267 => to_slv(opcode_type, 16#09#),
      268 => to_slv(opcode_type, 16#10#),
      269 => to_slv(opcode_type, 16#0D#),
      270 => to_slv(opcode_type, 16#05#),
      271 => to_slv(opcode_type, 16#04#),
      272 => to_slv(opcode_type, 16#0D#),
      273 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#06#),
      289 => to_slv(opcode_type, 16#06#),
      290 => to_slv(opcode_type, 16#01#),
      291 => to_slv(opcode_type, 16#09#),
      292 => to_slv(opcode_type, 16#0C#),
      293 => to_slv(opcode_type, 16#10#),
      294 => to_slv(opcode_type, 16#08#),
      295 => to_slv(opcode_type, 16#03#),
      296 => to_slv(opcode_type, 16#11#),
      297 => to_slv(opcode_type, 16#04#),
      298 => to_slv(opcode_type, 16#0D#),
      299 => to_slv(opcode_type, 16#08#),
      300 => to_slv(opcode_type, 16#03#),
      301 => to_slv(opcode_type, 16#08#),
      302 => to_slv(opcode_type, 16#87#),
      303 => to_slv(opcode_type, 16#A4#),
      304 => to_slv(opcode_type, 16#0E#),
      305 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#07#),
      321 => to_slv(opcode_type, 16#01#),
      322 => to_slv(opcode_type, 16#01#),
      323 => to_slv(opcode_type, 16#06#),
      324 => to_slv(opcode_type, 16#11#),
      325 => to_slv(opcode_type, 16#0F#),
      326 => to_slv(opcode_type, 16#08#),
      327 => to_slv(opcode_type, 16#03#),
      328 => to_slv(opcode_type, 16#07#),
      329 => to_slv(opcode_type, 16#0D#),
      330 => to_slv(opcode_type, 16#0A#),
      331 => to_slv(opcode_type, 16#09#),
      332 => to_slv(opcode_type, 16#06#),
      333 => to_slv(opcode_type, 16#11#),
      334 => to_slv(opcode_type, 16#0B#),
      335 => to_slv(opcode_type, 16#04#),
      336 => to_slv(opcode_type, 16#0C#),
      337 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#06#),
      353 => to_slv(opcode_type, 16#06#),
      354 => to_slv(opcode_type, 16#06#),
      355 => to_slv(opcode_type, 16#03#),
      356 => to_slv(opcode_type, 16#0D#),
      357 => to_slv(opcode_type, 16#02#),
      358 => to_slv(opcode_type, 16#10#),
      359 => to_slv(opcode_type, 16#09#),
      360 => to_slv(opcode_type, 16#09#),
      361 => to_slv(opcode_type, 16#0E#),
      362 => to_slv(opcode_type, 16#0F#),
      363 => to_slv(opcode_type, 16#04#),
      364 => to_slv(opcode_type, 16#0B#),
      365 => to_slv(opcode_type, 16#07#),
      366 => to_slv(opcode_type, 16#01#),
      367 => to_slv(opcode_type, 16#0A#),
      368 => to_slv(opcode_type, 16#10#),
      369 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#08#),
      385 => to_slv(opcode_type, 16#04#),
      386 => to_slv(opcode_type, 16#02#),
      387 => to_slv(opcode_type, 16#02#),
      388 => to_slv(opcode_type, 16#0F#),
      389 => to_slv(opcode_type, 16#07#),
      390 => to_slv(opcode_type, 16#02#),
      391 => to_slv(opcode_type, 16#06#),
      392 => to_slv(opcode_type, 16#0C#),
      393 => to_slv(opcode_type, 16#11#),
      394 => to_slv(opcode_type, 16#08#),
      395 => to_slv(opcode_type, 16#07#),
      396 => to_slv(opcode_type, 16#10#),
      397 => to_slv(opcode_type, 16#0D#),
      398 => to_slv(opcode_type, 16#08#),
      399 => to_slv(opcode_type, 16#11#),
      400 => to_slv(opcode_type, 16#10#),
      401 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#09#),
      417 => to_slv(opcode_type, 16#09#),
      418 => to_slv(opcode_type, 16#08#),
      419 => to_slv(opcode_type, 16#03#),
      420 => to_slv(opcode_type, 16#0D#),
      421 => to_slv(opcode_type, 16#05#),
      422 => to_slv(opcode_type, 16#0E#),
      423 => to_slv(opcode_type, 16#04#),
      424 => to_slv(opcode_type, 16#01#),
      425 => to_slv(opcode_type, 16#0B#),
      426 => to_slv(opcode_type, 16#05#),
      427 => to_slv(opcode_type, 16#07#),
      428 => to_slv(opcode_type, 16#03#),
      429 => to_slv(opcode_type, 16#0A#),
      430 => to_slv(opcode_type, 16#06#),
      431 => to_slv(opcode_type, 16#11#),
      432 => to_slv(opcode_type, 16#0D#),
      433 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#09#),
      449 => to_slv(opcode_type, 16#04#),
      450 => to_slv(opcode_type, 16#01#),
      451 => to_slv(opcode_type, 16#04#),
      452 => to_slv(opcode_type, 16#0B#),
      453 => to_slv(opcode_type, 16#08#),
      454 => to_slv(opcode_type, 16#05#),
      455 => to_slv(opcode_type, 16#06#),
      456 => to_slv(opcode_type, 16#0A#),
      457 => to_slv(opcode_type, 16#0A#),
      458 => to_slv(opcode_type, 16#08#),
      459 => to_slv(opcode_type, 16#07#),
      460 => to_slv(opcode_type, 16#10#),
      461 => to_slv(opcode_type, 16#0A#),
      462 => to_slv(opcode_type, 16#07#),
      463 => to_slv(opcode_type, 16#DF#),
      464 => to_slv(opcode_type, 16#0E#),
      465 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#07#),
      481 => to_slv(opcode_type, 16#04#),
      482 => to_slv(opcode_type, 16#09#),
      483 => to_slv(opcode_type, 16#03#),
      484 => to_slv(opcode_type, 16#0D#),
      485 => to_slv(opcode_type, 16#01#),
      486 => to_slv(opcode_type, 16#0E#),
      487 => to_slv(opcode_type, 16#07#),
      488 => to_slv(opcode_type, 16#03#),
      489 => to_slv(opcode_type, 16#09#),
      490 => to_slv(opcode_type, 16#10#),
      491 => to_slv(opcode_type, 16#0D#),
      492 => to_slv(opcode_type, 16#09#),
      493 => to_slv(opcode_type, 16#01#),
      494 => to_slv(opcode_type, 16#2A#),
      495 => to_slv(opcode_type, 16#05#),
      496 => to_slv(opcode_type, 16#0C#),
      497 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#05#),
      514 => to_slv(opcode_type, 16#09#),
      515 => to_slv(opcode_type, 16#06#),
      516 => to_slv(opcode_type, 16#10#),
      517 => to_slv(opcode_type, 16#0E#),
      518 => to_slv(opcode_type, 16#01#),
      519 => to_slv(opcode_type, 16#0B#),
      520 => to_slv(opcode_type, 16#08#),
      521 => to_slv(opcode_type, 16#02#),
      522 => to_slv(opcode_type, 16#04#),
      523 => to_slv(opcode_type, 16#0A#),
      524 => to_slv(opcode_type, 16#06#),
      525 => to_slv(opcode_type, 16#03#),
      526 => to_slv(opcode_type, 16#0D#),
      527 => to_slv(opcode_type, 16#01#),
      528 => to_slv(opcode_type, 16#3E#),
      529 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#09#),
      545 => to_slv(opcode_type, 16#05#),
      546 => to_slv(opcode_type, 16#05#),
      547 => to_slv(opcode_type, 16#06#),
      548 => to_slv(opcode_type, 16#0D#),
      549 => to_slv(opcode_type, 16#0F#),
      550 => to_slv(opcode_type, 16#08#),
      551 => to_slv(opcode_type, 16#04#),
      552 => to_slv(opcode_type, 16#04#),
      553 => to_slv(opcode_type, 16#0F#),
      554 => to_slv(opcode_type, 16#07#),
      555 => to_slv(opcode_type, 16#08#),
      556 => to_slv(opcode_type, 16#0A#),
      557 => to_slv(opcode_type, 16#88#),
      558 => to_slv(opcode_type, 16#09#),
      559 => to_slv(opcode_type, 16#0B#),
      560 => to_slv(opcode_type, 16#11#),
      561 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#09#),
      577 => to_slv(opcode_type, 16#08#),
      578 => to_slv(opcode_type, 16#06#),
      579 => to_slv(opcode_type, 16#08#),
      580 => to_slv(opcode_type, 16#86#),
      581 => to_slv(opcode_type, 16#11#),
      582 => to_slv(opcode_type, 16#05#),
      583 => to_slv(opcode_type, 16#11#),
      584 => to_slv(opcode_type, 16#02#),
      585 => to_slv(opcode_type, 16#09#),
      586 => to_slv(opcode_type, 16#0B#),
      587 => to_slv(opcode_type, 16#0B#),
      588 => to_slv(opcode_type, 16#09#),
      589 => to_slv(opcode_type, 16#07#),
      590 => to_slv(opcode_type, 16#10#),
      591 => to_slv(opcode_type, 16#9B#),
      592 => to_slv(opcode_type, 16#0E#),
      593 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#08#),
      609 => to_slv(opcode_type, 16#04#),
      610 => to_slv(opcode_type, 16#04#),
      611 => to_slv(opcode_type, 16#01#),
      612 => to_slv(opcode_type, 16#0C#),
      613 => to_slv(opcode_type, 16#06#),
      614 => to_slv(opcode_type, 16#08#),
      615 => to_slv(opcode_type, 16#08#),
      616 => to_slv(opcode_type, 16#11#),
      617 => to_slv(opcode_type, 16#10#),
      618 => to_slv(opcode_type, 16#01#),
      619 => to_slv(opcode_type, 16#0B#),
      620 => to_slv(opcode_type, 16#09#),
      621 => to_slv(opcode_type, 16#01#),
      622 => to_slv(opcode_type, 16#11#),
      623 => to_slv(opcode_type, 16#04#),
      624 => to_slv(opcode_type, 16#0E#),
      625 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#09#),
      641 => to_slv(opcode_type, 16#03#),
      642 => to_slv(opcode_type, 16#07#),
      643 => to_slv(opcode_type, 16#07#),
      644 => to_slv(opcode_type, 16#0E#),
      645 => to_slv(opcode_type, 16#0E#),
      646 => to_slv(opcode_type, 16#08#),
      647 => to_slv(opcode_type, 16#92#),
      648 => to_slv(opcode_type, 16#11#),
      649 => to_slv(opcode_type, 16#03#),
      650 => to_slv(opcode_type, 16#08#),
      651 => to_slv(opcode_type, 16#07#),
      652 => to_slv(opcode_type, 16#0B#),
      653 => to_slv(opcode_type, 16#E2#),
      654 => to_slv(opcode_type, 16#07#),
      655 => to_slv(opcode_type, 16#11#),
      656 => to_slv(opcode_type, 16#0D#),
      657 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#07#),
      673 => to_slv(opcode_type, 16#04#),
      674 => to_slv(opcode_type, 16#03#),
      675 => to_slv(opcode_type, 16#03#),
      676 => to_slv(opcode_type, 16#54#),
      677 => to_slv(opcode_type, 16#06#),
      678 => to_slv(opcode_type, 16#06#),
      679 => to_slv(opcode_type, 16#01#),
      680 => to_slv(opcode_type, 16#0B#),
      681 => to_slv(opcode_type, 16#08#),
      682 => to_slv(opcode_type, 16#0C#),
      683 => to_slv(opcode_type, 16#0D#),
      684 => to_slv(opcode_type, 16#07#),
      685 => to_slv(opcode_type, 16#05#),
      686 => to_slv(opcode_type, 16#0D#),
      687 => to_slv(opcode_type, 16#01#),
      688 => to_slv(opcode_type, 16#11#),
      689 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#06#),
      705 => to_slv(opcode_type, 16#01#),
      706 => to_slv(opcode_type, 16#05#),
      707 => to_slv(opcode_type, 16#06#),
      708 => to_slv(opcode_type, 16#11#),
      709 => to_slv(opcode_type, 16#0F#),
      710 => to_slv(opcode_type, 16#07#),
      711 => to_slv(opcode_type, 16#01#),
      712 => to_slv(opcode_type, 16#04#),
      713 => to_slv(opcode_type, 16#1D#),
      714 => to_slv(opcode_type, 16#07#),
      715 => to_slv(opcode_type, 16#07#),
      716 => to_slv(opcode_type, 16#0C#),
      717 => to_slv(opcode_type, 16#0E#),
      718 => to_slv(opcode_type, 16#06#),
      719 => to_slv(opcode_type, 16#6E#),
      720 => to_slv(opcode_type, 16#BC#),
      721 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#07#),
      737 => to_slv(opcode_type, 16#03#),
      738 => to_slv(opcode_type, 16#06#),
      739 => to_slv(opcode_type, 16#04#),
      740 => to_slv(opcode_type, 16#0E#),
      741 => to_slv(opcode_type, 16#04#),
      742 => to_slv(opcode_type, 16#11#),
      743 => to_slv(opcode_type, 16#06#),
      744 => to_slv(opcode_type, 16#09#),
      745 => to_slv(opcode_type, 16#05#),
      746 => to_slv(opcode_type, 16#0A#),
      747 => to_slv(opcode_type, 16#05#),
      748 => to_slv(opcode_type, 16#0B#),
      749 => to_slv(opcode_type, 16#06#),
      750 => to_slv(opcode_type, 16#01#),
      751 => to_slv(opcode_type, 16#0A#),
      752 => to_slv(opcode_type, 16#0D#),
      753 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#09#),
      769 => to_slv(opcode_type, 16#05#),
      770 => to_slv(opcode_type, 16#02#),
      771 => to_slv(opcode_type, 16#03#),
      772 => to_slv(opcode_type, 16#0C#),
      773 => to_slv(opcode_type, 16#07#),
      774 => to_slv(opcode_type, 16#02#),
      775 => to_slv(opcode_type, 16#07#),
      776 => to_slv(opcode_type, 16#0A#),
      777 => to_slv(opcode_type, 16#0E#),
      778 => to_slv(opcode_type, 16#07#),
      779 => to_slv(opcode_type, 16#07#),
      780 => to_slv(opcode_type, 16#11#),
      781 => to_slv(opcode_type, 16#0B#),
      782 => to_slv(opcode_type, 16#09#),
      783 => to_slv(opcode_type, 16#11#),
      784 => to_slv(opcode_type, 16#0B#),
      785 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#08#),
      801 => to_slv(opcode_type, 16#04#),
      802 => to_slv(opcode_type, 16#09#),
      803 => to_slv(opcode_type, 16#02#),
      804 => to_slv(opcode_type, 16#D9#),
      805 => to_slv(opcode_type, 16#02#),
      806 => to_slv(opcode_type, 16#10#),
      807 => to_slv(opcode_type, 16#06#),
      808 => to_slv(opcode_type, 16#07#),
      809 => to_slv(opcode_type, 16#01#),
      810 => to_slv(opcode_type, 16#10#),
      811 => to_slv(opcode_type, 16#08#),
      812 => to_slv(opcode_type, 16#0A#),
      813 => to_slv(opcode_type, 16#EF#),
      814 => to_slv(opcode_type, 16#05#),
      815 => to_slv(opcode_type, 16#05#),
      816 => to_slv(opcode_type, 16#0E#),
      817 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#09#),
      833 => to_slv(opcode_type, 16#09#),
      834 => to_slv(opcode_type, 16#08#),
      835 => to_slv(opcode_type, 16#06#),
      836 => to_slv(opcode_type, 16#0B#),
      837 => to_slv(opcode_type, 16#0B#),
      838 => to_slv(opcode_type, 16#07#),
      839 => to_slv(opcode_type, 16#10#),
      840 => to_slv(opcode_type, 16#22#),
      841 => to_slv(opcode_type, 16#08#),
      842 => to_slv(opcode_type, 16#08#),
      843 => to_slv(opcode_type, 16#0F#),
      844 => to_slv(opcode_type, 16#0C#),
      845 => to_slv(opcode_type, 16#01#),
      846 => to_slv(opcode_type, 16#11#),
      847 => to_slv(opcode_type, 16#03#),
      848 => to_slv(opcode_type, 16#76#),
      849 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#07#),
      865 => to_slv(opcode_type, 16#06#),
      866 => to_slv(opcode_type, 16#05#),
      867 => to_slv(opcode_type, 16#01#),
      868 => to_slv(opcode_type, 16#11#),
      869 => to_slv(opcode_type, 16#04#),
      870 => to_slv(opcode_type, 16#07#),
      871 => to_slv(opcode_type, 16#0E#),
      872 => to_slv(opcode_type, 16#0C#),
      873 => to_slv(opcode_type, 16#07#),
      874 => to_slv(opcode_type, 16#01#),
      875 => to_slv(opcode_type, 16#01#),
      876 => to_slv(opcode_type, 16#0A#),
      877 => to_slv(opcode_type, 16#01#),
      878 => to_slv(opcode_type, 16#09#),
      879 => to_slv(opcode_type, 16#11#),
      880 => to_slv(opcode_type, 16#10#),
      881 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#08#),
      898 => to_slv(opcode_type, 16#09#),
      899 => to_slv(opcode_type, 16#09#),
      900 => to_slv(opcode_type, 16#0B#),
      901 => to_slv(opcode_type, 16#0B#),
      902 => to_slv(opcode_type, 16#09#),
      903 => to_slv(opcode_type, 16#0C#),
      904 => to_slv(opcode_type, 16#0B#),
      905 => to_slv(opcode_type, 16#03#),
      906 => to_slv(opcode_type, 16#03#),
      907 => to_slv(opcode_type, 16#0D#),
      908 => to_slv(opcode_type, 16#01#),
      909 => to_slv(opcode_type, 16#04#),
      910 => to_slv(opcode_type, 16#08#),
      911 => to_slv(opcode_type, 16#0A#),
      912 => to_slv(opcode_type, 16#10#),
      913 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#08#),
      929 => to_slv(opcode_type, 16#09#),
      930 => to_slv(opcode_type, 16#03#),
      931 => to_slv(opcode_type, 16#03#),
      932 => to_slv(opcode_type, 16#0C#),
      933 => to_slv(opcode_type, 16#03#),
      934 => to_slv(opcode_type, 16#06#),
      935 => to_slv(opcode_type, 16#1E#),
      936 => to_slv(opcode_type, 16#10#),
      937 => to_slv(opcode_type, 16#05#),
      938 => to_slv(opcode_type, 16#07#),
      939 => to_slv(opcode_type, 16#09#),
      940 => to_slv(opcode_type, 16#10#),
      941 => to_slv(opcode_type, 16#0B#),
      942 => to_slv(opcode_type, 16#09#),
      943 => to_slv(opcode_type, 16#0F#),
      944 => to_slv(opcode_type, 16#1A#),
      945 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#01#),
      962 => to_slv(opcode_type, 16#06#),
      963 => to_slv(opcode_type, 16#06#),
      964 => to_slv(opcode_type, 16#CF#),
      965 => to_slv(opcode_type, 16#0F#),
      966 => to_slv(opcode_type, 16#06#),
      967 => to_slv(opcode_type, 16#0D#),
      968 => to_slv(opcode_type, 16#0C#),
      969 => to_slv(opcode_type, 16#02#),
      970 => to_slv(opcode_type, 16#06#),
      971 => to_slv(opcode_type, 16#09#),
      972 => to_slv(opcode_type, 16#0F#),
      973 => to_slv(opcode_type, 16#0D#),
      974 => to_slv(opcode_type, 16#07#),
      975 => to_slv(opcode_type, 16#0D#),
      976 => to_slv(opcode_type, 16#0C#),
      977 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#06#),
      993 => to_slv(opcode_type, 16#08#),
      994 => to_slv(opcode_type, 16#04#),
      995 => to_slv(opcode_type, 16#09#),
      996 => to_slv(opcode_type, 16#80#),
      997 => to_slv(opcode_type, 16#0F#),
      998 => to_slv(opcode_type, 16#03#),
      999 => to_slv(opcode_type, 16#04#),
      1000 => to_slv(opcode_type, 16#0D#),
      1001 => to_slv(opcode_type, 16#09#),
      1002 => to_slv(opcode_type, 16#07#),
      1003 => to_slv(opcode_type, 16#02#),
      1004 => to_slv(opcode_type, 16#0E#),
      1005 => to_slv(opcode_type, 16#09#),
      1006 => to_slv(opcode_type, 16#6F#),
      1007 => to_slv(opcode_type, 16#0B#),
      1008 => to_slv(opcode_type, 16#0F#),
      1009 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#07#),
      1025 => to_slv(opcode_type, 16#08#),
      1026 => to_slv(opcode_type, 16#01#),
      1027 => to_slv(opcode_type, 16#03#),
      1028 => to_slv(opcode_type, 16#0B#),
      1029 => to_slv(opcode_type, 16#09#),
      1030 => to_slv(opcode_type, 16#08#),
      1031 => to_slv(opcode_type, 16#0B#),
      1032 => to_slv(opcode_type, 16#11#),
      1033 => to_slv(opcode_type, 16#03#),
      1034 => to_slv(opcode_type, 16#0A#),
      1035 => to_slv(opcode_type, 16#03#),
      1036 => to_slv(opcode_type, 16#07#),
      1037 => to_slv(opcode_type, 16#03#),
      1038 => to_slv(opcode_type, 16#11#),
      1039 => to_slv(opcode_type, 16#03#),
      1040 => to_slv(opcode_type, 16#0D#),
      1041 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#06#),
      1057 => to_slv(opcode_type, 16#06#),
      1058 => to_slv(opcode_type, 16#09#),
      1059 => to_slv(opcode_type, 16#01#),
      1060 => to_slv(opcode_type, 16#0B#),
      1061 => to_slv(opcode_type, 16#02#),
      1062 => to_slv(opcode_type, 16#10#),
      1063 => to_slv(opcode_type, 16#03#),
      1064 => to_slv(opcode_type, 16#05#),
      1065 => to_slv(opcode_type, 16#10#),
      1066 => to_slv(opcode_type, 16#01#),
      1067 => to_slv(opcode_type, 16#07#),
      1068 => to_slv(opcode_type, 16#09#),
      1069 => to_slv(opcode_type, 16#0D#),
      1070 => to_slv(opcode_type, 16#0C#),
      1071 => to_slv(opcode_type, 16#05#),
      1072 => to_slv(opcode_type, 16#11#),
      1073 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#09#),
      1089 => to_slv(opcode_type, 16#03#),
      1090 => to_slv(opcode_type, 16#09#),
      1091 => to_slv(opcode_type, 16#04#),
      1092 => to_slv(opcode_type, 16#11#),
      1093 => to_slv(opcode_type, 16#01#),
      1094 => to_slv(opcode_type, 16#0D#),
      1095 => to_slv(opcode_type, 16#08#),
      1096 => to_slv(opcode_type, 16#02#),
      1097 => to_slv(opcode_type, 16#04#),
      1098 => to_slv(opcode_type, 16#0F#),
      1099 => to_slv(opcode_type, 16#08#),
      1100 => to_slv(opcode_type, 16#02#),
      1101 => to_slv(opcode_type, 16#10#),
      1102 => to_slv(opcode_type, 16#09#),
      1103 => to_slv(opcode_type, 16#0A#),
      1104 => to_slv(opcode_type, 16#0C#),
      1105 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#06#),
      1121 => to_slv(opcode_type, 16#06#),
      1122 => to_slv(opcode_type, 16#06#),
      1123 => to_slv(opcode_type, 16#09#),
      1124 => to_slv(opcode_type, 16#0F#),
      1125 => to_slv(opcode_type, 16#10#),
      1126 => to_slv(opcode_type, 16#09#),
      1127 => to_slv(opcode_type, 16#0F#),
      1128 => to_slv(opcode_type, 16#0E#),
      1129 => to_slv(opcode_type, 16#07#),
      1130 => to_slv(opcode_type, 16#05#),
      1131 => to_slv(opcode_type, 16#0B#),
      1132 => to_slv(opcode_type, 16#04#),
      1133 => to_slv(opcode_type, 16#10#),
      1134 => to_slv(opcode_type, 16#01#),
      1135 => to_slv(opcode_type, 16#01#),
      1136 => to_slv(opcode_type, 16#0F#),
      1137 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#06#),
      1153 => to_slv(opcode_type, 16#03#),
      1154 => to_slv(opcode_type, 16#01#),
      1155 => to_slv(opcode_type, 16#04#),
      1156 => to_slv(opcode_type, 16#0E#),
      1157 => to_slv(opcode_type, 16#07#),
      1158 => to_slv(opcode_type, 16#04#),
      1159 => to_slv(opcode_type, 16#07#),
      1160 => to_slv(opcode_type, 16#0F#),
      1161 => to_slv(opcode_type, 16#0A#),
      1162 => to_slv(opcode_type, 16#07#),
      1163 => to_slv(opcode_type, 16#07#),
      1164 => to_slv(opcode_type, 16#0A#),
      1165 => to_slv(opcode_type, 16#10#),
      1166 => to_slv(opcode_type, 16#07#),
      1167 => to_slv(opcode_type, 16#13#),
      1168 => to_slv(opcode_type, 16#10#),
      1169 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#08#),
      1185 => to_slv(opcode_type, 16#02#),
      1186 => to_slv(opcode_type, 16#06#),
      1187 => to_slv(opcode_type, 16#07#),
      1188 => to_slv(opcode_type, 16#0C#),
      1189 => to_slv(opcode_type, 16#0E#),
      1190 => to_slv(opcode_type, 16#07#),
      1191 => to_slv(opcode_type, 16#0A#),
      1192 => to_slv(opcode_type, 16#7E#),
      1193 => to_slv(opcode_type, 16#08#),
      1194 => to_slv(opcode_type, 16#05#),
      1195 => to_slv(opcode_type, 16#07#),
      1196 => to_slv(opcode_type, 16#0E#),
      1197 => to_slv(opcode_type, 16#18#),
      1198 => to_slv(opcode_type, 16#06#),
      1199 => to_slv(opcode_type, 16#0A#),
      1200 => to_slv(opcode_type, 16#0E#),
      1201 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#06#),
      1217 => to_slv(opcode_type, 16#05#),
      1218 => to_slv(opcode_type, 16#05#),
      1219 => to_slv(opcode_type, 16#07#),
      1220 => to_slv(opcode_type, 16#7E#),
      1221 => to_slv(opcode_type, 16#10#),
      1222 => to_slv(opcode_type, 16#09#),
      1223 => to_slv(opcode_type, 16#09#),
      1224 => to_slv(opcode_type, 16#04#),
      1225 => to_slv(opcode_type, 16#0C#),
      1226 => to_slv(opcode_type, 16#08#),
      1227 => to_slv(opcode_type, 16#3A#),
      1228 => to_slv(opcode_type, 16#0B#),
      1229 => to_slv(opcode_type, 16#04#),
      1230 => to_slv(opcode_type, 16#08#),
      1231 => to_slv(opcode_type, 16#0E#),
      1232 => to_slv(opcode_type, 16#10#),
      1233 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#09#),
      1249 => to_slv(opcode_type, 16#02#),
      1250 => to_slv(opcode_type, 16#08#),
      1251 => to_slv(opcode_type, 16#04#),
      1252 => to_slv(opcode_type, 16#0D#),
      1253 => to_slv(opcode_type, 16#01#),
      1254 => to_slv(opcode_type, 16#0C#),
      1255 => to_slv(opcode_type, 16#08#),
      1256 => to_slv(opcode_type, 16#09#),
      1257 => to_slv(opcode_type, 16#08#),
      1258 => to_slv(opcode_type, 16#0A#),
      1259 => to_slv(opcode_type, 16#11#),
      1260 => to_slv(opcode_type, 16#04#),
      1261 => to_slv(opcode_type, 16#0F#),
      1262 => to_slv(opcode_type, 16#08#),
      1263 => to_slv(opcode_type, 16#0F#),
      1264 => to_slv(opcode_type, 16#0A#),
      1265 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#04#),
      1282 => to_slv(opcode_type, 16#02#),
      1283 => to_slv(opcode_type, 16#06#),
      1284 => to_slv(opcode_type, 16#10#),
      1285 => to_slv(opcode_type, 16#11#),
      1286 => to_slv(opcode_type, 16#06#),
      1287 => to_slv(opcode_type, 16#02#),
      1288 => to_slv(opcode_type, 16#01#),
      1289 => to_slv(opcode_type, 16#0D#),
      1290 => to_slv(opcode_type, 16#09#),
      1291 => to_slv(opcode_type, 16#07#),
      1292 => to_slv(opcode_type, 16#0F#),
      1293 => to_slv(opcode_type, 16#0C#),
      1294 => to_slv(opcode_type, 16#08#),
      1295 => to_slv(opcode_type, 16#0A#),
      1296 => to_slv(opcode_type, 16#0F#),
      1297 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#06#),
      1313 => to_slv(opcode_type, 16#01#),
      1314 => to_slv(opcode_type, 16#01#),
      1315 => to_slv(opcode_type, 16#04#),
      1316 => to_slv(opcode_type, 16#0B#),
      1317 => to_slv(opcode_type, 16#06#),
      1318 => to_slv(opcode_type, 16#06#),
      1319 => to_slv(opcode_type, 16#01#),
      1320 => to_slv(opcode_type, 16#0B#),
      1321 => to_slv(opcode_type, 16#05#),
      1322 => to_slv(opcode_type, 16#0A#),
      1323 => to_slv(opcode_type, 16#08#),
      1324 => to_slv(opcode_type, 16#04#),
      1325 => to_slv(opcode_type, 16#0B#),
      1326 => to_slv(opcode_type, 16#08#),
      1327 => to_slv(opcode_type, 16#10#),
      1328 => to_slv(opcode_type, 16#11#),
      1329 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#07#),
      1345 => to_slv(opcode_type, 16#07#),
      1346 => to_slv(opcode_type, 16#07#),
      1347 => to_slv(opcode_type, 16#03#),
      1348 => to_slv(opcode_type, 16#92#),
      1349 => to_slv(opcode_type, 16#08#),
      1350 => to_slv(opcode_type, 16#0B#),
      1351 => to_slv(opcode_type, 16#0E#),
      1352 => to_slv(opcode_type, 16#01#),
      1353 => to_slv(opcode_type, 16#04#),
      1354 => to_slv(opcode_type, 16#10#),
      1355 => to_slv(opcode_type, 16#04#),
      1356 => to_slv(opcode_type, 16#07#),
      1357 => to_slv(opcode_type, 16#05#),
      1358 => to_slv(opcode_type, 16#0A#),
      1359 => to_slv(opcode_type, 16#01#),
      1360 => to_slv(opcode_type, 16#0B#),
      1361 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#09#),
      1377 => to_slv(opcode_type, 16#06#),
      1378 => to_slv(opcode_type, 16#08#),
      1379 => to_slv(opcode_type, 16#03#),
      1380 => to_slv(opcode_type, 16#0D#),
      1381 => to_slv(opcode_type, 16#09#),
      1382 => to_slv(opcode_type, 16#DD#),
      1383 => to_slv(opcode_type, 16#1E#),
      1384 => to_slv(opcode_type, 16#05#),
      1385 => to_slv(opcode_type, 16#09#),
      1386 => to_slv(opcode_type, 16#0F#),
      1387 => to_slv(opcode_type, 16#26#),
      1388 => to_slv(opcode_type, 16#02#),
      1389 => to_slv(opcode_type, 16#08#),
      1390 => to_slv(opcode_type, 16#01#),
      1391 => to_slv(opcode_type, 16#19#),
      1392 => to_slv(opcode_type, 16#0F#),
      1393 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#07#),
      1410 => to_slv(opcode_type, 16#05#),
      1411 => to_slv(opcode_type, 16#03#),
      1412 => to_slv(opcode_type, 16#0E#),
      1413 => to_slv(opcode_type, 16#02#),
      1414 => to_slv(opcode_type, 16#04#),
      1415 => to_slv(opcode_type, 16#A4#),
      1416 => to_slv(opcode_type, 16#08#),
      1417 => to_slv(opcode_type, 16#08#),
      1418 => to_slv(opcode_type, 16#08#),
      1419 => to_slv(opcode_type, 16#AA#),
      1420 => to_slv(opcode_type, 16#0F#),
      1421 => to_slv(opcode_type, 16#02#),
      1422 => to_slv(opcode_type, 16#0D#),
      1423 => to_slv(opcode_type, 16#05#),
      1424 => to_slv(opcode_type, 16#0A#),
      1425 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#06#),
      1441 => to_slv(opcode_type, 16#03#),
      1442 => to_slv(opcode_type, 16#09#),
      1443 => to_slv(opcode_type, 16#06#),
      1444 => to_slv(opcode_type, 16#0D#),
      1445 => to_slv(opcode_type, 16#0B#),
      1446 => to_slv(opcode_type, 16#02#),
      1447 => to_slv(opcode_type, 16#0C#),
      1448 => to_slv(opcode_type, 16#06#),
      1449 => to_slv(opcode_type, 16#08#),
      1450 => to_slv(opcode_type, 16#07#),
      1451 => to_slv(opcode_type, 16#0D#),
      1452 => to_slv(opcode_type, 16#0A#),
      1453 => to_slv(opcode_type, 16#03#),
      1454 => to_slv(opcode_type, 16#85#),
      1455 => to_slv(opcode_type, 16#04#),
      1456 => to_slv(opcode_type, 16#FE#),
      1457 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#09#),
      1473 => to_slv(opcode_type, 16#05#),
      1474 => to_slv(opcode_type, 16#05#),
      1475 => to_slv(opcode_type, 16#08#),
      1476 => to_slv(opcode_type, 16#0B#),
      1477 => to_slv(opcode_type, 16#0D#),
      1478 => to_slv(opcode_type, 16#06#),
      1479 => to_slv(opcode_type, 16#09#),
      1480 => to_slv(opcode_type, 16#09#),
      1481 => to_slv(opcode_type, 16#0C#),
      1482 => to_slv(opcode_type, 16#10#),
      1483 => to_slv(opcode_type, 16#07#),
      1484 => to_slv(opcode_type, 16#0B#),
      1485 => to_slv(opcode_type, 16#10#),
      1486 => to_slv(opcode_type, 16#05#),
      1487 => to_slv(opcode_type, 16#04#),
      1488 => to_slv(opcode_type, 16#0C#),
      1489 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#07#),
      1505 => to_slv(opcode_type, 16#05#),
      1506 => to_slv(opcode_type, 16#03#),
      1507 => to_slv(opcode_type, 16#07#),
      1508 => to_slv(opcode_type, 16#10#),
      1509 => to_slv(opcode_type, 16#0D#),
      1510 => to_slv(opcode_type, 16#06#),
      1511 => to_slv(opcode_type, 16#09#),
      1512 => to_slv(opcode_type, 16#05#),
      1513 => to_slv(opcode_type, 16#0E#),
      1514 => to_slv(opcode_type, 16#07#),
      1515 => to_slv(opcode_type, 16#0D#),
      1516 => to_slv(opcode_type, 16#0E#),
      1517 => to_slv(opcode_type, 16#02#),
      1518 => to_slv(opcode_type, 16#06#),
      1519 => to_slv(opcode_type, 16#11#),
      1520 => to_slv(opcode_type, 16#0C#),
      1521 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#07#),
      1537 => to_slv(opcode_type, 16#03#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#04#),
      1540 => to_slv(opcode_type, 16#0F#),
      1541 => to_slv(opcode_type, 16#04#),
      1542 => to_slv(opcode_type, 16#0E#),
      1543 => to_slv(opcode_type, 16#07#),
      1544 => to_slv(opcode_type, 16#09#),
      1545 => to_slv(opcode_type, 16#06#),
      1546 => to_slv(opcode_type, 16#0E#),
      1547 => to_slv(opcode_type, 16#10#),
      1548 => to_slv(opcode_type, 16#04#),
      1549 => to_slv(opcode_type, 16#0E#),
      1550 => to_slv(opcode_type, 16#07#),
      1551 => to_slv(opcode_type, 16#0E#),
      1552 => to_slv(opcode_type, 16#0A#),
      1553 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#09#),
      1569 => to_slv(opcode_type, 16#07#),
      1570 => to_slv(opcode_type, 16#04#),
      1571 => to_slv(opcode_type, 16#09#),
      1572 => to_slv(opcode_type, 16#15#),
      1573 => to_slv(opcode_type, 16#0E#),
      1574 => to_slv(opcode_type, 16#07#),
      1575 => to_slv(opcode_type, 16#03#),
      1576 => to_slv(opcode_type, 16#0C#),
      1577 => to_slv(opcode_type, 16#09#),
      1578 => to_slv(opcode_type, 16#10#),
      1579 => to_slv(opcode_type, 16#67#),
      1580 => to_slv(opcode_type, 16#06#),
      1581 => to_slv(opcode_type, 16#07#),
      1582 => to_slv(opcode_type, 16#0A#),
      1583 => to_slv(opcode_type, 16#0E#),
      1584 => to_slv(opcode_type, 16#A1#),
      1585 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#08#),
      1601 => to_slv(opcode_type, 16#01#),
      1602 => to_slv(opcode_type, 16#03#),
      1603 => to_slv(opcode_type, 16#06#),
      1604 => to_slv(opcode_type, 16#10#),
      1605 => to_slv(opcode_type, 16#10#),
      1606 => to_slv(opcode_type, 16#08#),
      1607 => to_slv(opcode_type, 16#01#),
      1608 => to_slv(opcode_type, 16#02#),
      1609 => to_slv(opcode_type, 16#0A#),
      1610 => to_slv(opcode_type, 16#08#),
      1611 => to_slv(opcode_type, 16#08#),
      1612 => to_slv(opcode_type, 16#11#),
      1613 => to_slv(opcode_type, 16#0C#),
      1614 => to_slv(opcode_type, 16#06#),
      1615 => to_slv(opcode_type, 16#0B#),
      1616 => to_slv(opcode_type, 16#0E#),
      1617 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#06#),
      1633 => to_slv(opcode_type, 16#08#),
      1634 => to_slv(opcode_type, 16#02#),
      1635 => to_slv(opcode_type, 16#03#),
      1636 => to_slv(opcode_type, 16#0E#),
      1637 => to_slv(opcode_type, 16#03#),
      1638 => to_slv(opcode_type, 16#03#),
      1639 => to_slv(opcode_type, 16#0F#),
      1640 => to_slv(opcode_type, 16#06#),
      1641 => to_slv(opcode_type, 16#07#),
      1642 => to_slv(opcode_type, 16#06#),
      1643 => to_slv(opcode_type, 16#0B#),
      1644 => to_slv(opcode_type, 16#0B#),
      1645 => to_slv(opcode_type, 16#08#),
      1646 => to_slv(opcode_type, 16#0E#),
      1647 => to_slv(opcode_type, 16#0A#),
      1648 => to_slv(opcode_type, 16#0E#),
      1649 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#03#),
      1666 => to_slv(opcode_type, 16#07#),
      1667 => to_slv(opcode_type, 16#09#),
      1668 => to_slv(opcode_type, 16#D4#),
      1669 => to_slv(opcode_type, 16#0F#),
      1670 => to_slv(opcode_type, 16#04#),
      1671 => to_slv(opcode_type, 16#0B#),
      1672 => to_slv(opcode_type, 16#09#),
      1673 => to_slv(opcode_type, 16#07#),
      1674 => to_slv(opcode_type, 16#04#),
      1675 => to_slv(opcode_type, 16#0B#),
      1676 => to_slv(opcode_type, 16#06#),
      1677 => to_slv(opcode_type, 16#0B#),
      1678 => to_slv(opcode_type, 16#91#),
      1679 => to_slv(opcode_type, 16#05#),
      1680 => to_slv(opcode_type, 16#0D#),
      1681 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#07#),
      1697 => to_slv(opcode_type, 16#01#),
      1698 => to_slv(opcode_type, 16#01#),
      1699 => to_slv(opcode_type, 16#06#),
      1700 => to_slv(opcode_type, 16#0E#),
      1701 => to_slv(opcode_type, 16#0C#),
      1702 => to_slv(opcode_type, 16#09#),
      1703 => to_slv(opcode_type, 16#01#),
      1704 => to_slv(opcode_type, 16#06#),
      1705 => to_slv(opcode_type, 16#0D#),
      1706 => to_slv(opcode_type, 16#11#),
      1707 => to_slv(opcode_type, 16#09#),
      1708 => to_slv(opcode_type, 16#03#),
      1709 => to_slv(opcode_type, 16#0F#),
      1710 => to_slv(opcode_type, 16#06#),
      1711 => to_slv(opcode_type, 16#39#),
      1712 => to_slv(opcode_type, 16#0A#),
      1713 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#08#),
      1729 => to_slv(opcode_type, 16#02#),
      1730 => to_slv(opcode_type, 16#07#),
      1731 => to_slv(opcode_type, 16#07#),
      1732 => to_slv(opcode_type, 16#0B#),
      1733 => to_slv(opcode_type, 16#10#),
      1734 => to_slv(opcode_type, 16#09#),
      1735 => to_slv(opcode_type, 16#0D#),
      1736 => to_slv(opcode_type, 16#50#),
      1737 => to_slv(opcode_type, 16#03#),
      1738 => to_slv(opcode_type, 16#08#),
      1739 => to_slv(opcode_type, 16#07#),
      1740 => to_slv(opcode_type, 16#0F#),
      1741 => to_slv(opcode_type, 16#0D#),
      1742 => to_slv(opcode_type, 16#08#),
      1743 => to_slv(opcode_type, 16#0A#),
      1744 => to_slv(opcode_type, 16#0F#),
      1745 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#09#),
      1761 => to_slv(opcode_type, 16#02#),
      1762 => to_slv(opcode_type, 16#04#),
      1763 => to_slv(opcode_type, 16#08#),
      1764 => to_slv(opcode_type, 16#11#),
      1765 => to_slv(opcode_type, 16#11#),
      1766 => to_slv(opcode_type, 16#06#),
      1767 => to_slv(opcode_type, 16#08#),
      1768 => to_slv(opcode_type, 16#08#),
      1769 => to_slv(opcode_type, 16#0F#),
      1770 => to_slv(opcode_type, 16#0D#),
      1771 => to_slv(opcode_type, 16#06#),
      1772 => to_slv(opcode_type, 16#0D#),
      1773 => to_slv(opcode_type, 16#F5#),
      1774 => to_slv(opcode_type, 16#02#),
      1775 => to_slv(opcode_type, 16#03#),
      1776 => to_slv(opcode_type, 16#0E#),
      1777 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#07#),
      1793 => to_slv(opcode_type, 16#09#),
      1794 => to_slv(opcode_type, 16#03#),
      1795 => to_slv(opcode_type, 16#01#),
      1796 => to_slv(opcode_type, 16#0E#),
      1797 => to_slv(opcode_type, 16#02#),
      1798 => to_slv(opcode_type, 16#08#),
      1799 => to_slv(opcode_type, 16#10#),
      1800 => to_slv(opcode_type, 16#5A#),
      1801 => to_slv(opcode_type, 16#01#),
      1802 => to_slv(opcode_type, 16#09#),
      1803 => to_slv(opcode_type, 16#08#),
      1804 => to_slv(opcode_type, 16#0C#),
      1805 => to_slv(opcode_type, 16#0F#),
      1806 => to_slv(opcode_type, 16#09#),
      1807 => to_slv(opcode_type, 16#0D#),
      1808 => to_slv(opcode_type, 16#0D#),
      1809 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#09#),
      1825 => to_slv(opcode_type, 16#01#),
      1826 => to_slv(opcode_type, 16#08#),
      1827 => to_slv(opcode_type, 16#02#),
      1828 => to_slv(opcode_type, 16#11#),
      1829 => to_slv(opcode_type, 16#06#),
      1830 => to_slv(opcode_type, 16#0A#),
      1831 => to_slv(opcode_type, 16#11#),
      1832 => to_slv(opcode_type, 16#08#),
      1833 => to_slv(opcode_type, 16#09#),
      1834 => to_slv(opcode_type, 16#02#),
      1835 => to_slv(opcode_type, 16#0D#),
      1836 => to_slv(opcode_type, 16#04#),
      1837 => to_slv(opcode_type, 16#10#),
      1838 => to_slv(opcode_type, 16#08#),
      1839 => to_slv(opcode_type, 16#0F#),
      1840 => to_slv(opcode_type, 16#0F#),
      1841 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#07#),
      1857 => to_slv(opcode_type, 16#08#),
      1858 => to_slv(opcode_type, 16#08#),
      1859 => to_slv(opcode_type, 16#07#),
      1860 => to_slv(opcode_type, 16#0C#),
      1861 => to_slv(opcode_type, 16#D8#),
      1862 => to_slv(opcode_type, 16#03#),
      1863 => to_slv(opcode_type, 16#11#),
      1864 => to_slv(opcode_type, 16#09#),
      1865 => to_slv(opcode_type, 16#01#),
      1866 => to_slv(opcode_type, 16#0F#),
      1867 => to_slv(opcode_type, 16#05#),
      1868 => to_slv(opcode_type, 16#0E#),
      1869 => to_slv(opcode_type, 16#06#),
      1870 => to_slv(opcode_type, 16#02#),
      1871 => to_slv(opcode_type, 16#11#),
      1872 => to_slv(opcode_type, 16#0B#),
      1873 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#08#),
      1890 => to_slv(opcode_type, 16#03#),
      1891 => to_slv(opcode_type, 16#05#),
      1892 => to_slv(opcode_type, 16#0C#),
      1893 => to_slv(opcode_type, 16#04#),
      1894 => to_slv(opcode_type, 16#03#),
      1895 => to_slv(opcode_type, 16#BA#),
      1896 => to_slv(opcode_type, 16#08#),
      1897 => to_slv(opcode_type, 16#03#),
      1898 => to_slv(opcode_type, 16#07#),
      1899 => to_slv(opcode_type, 16#0B#),
      1900 => to_slv(opcode_type, 16#0F#),
      1901 => to_slv(opcode_type, 16#09#),
      1902 => to_slv(opcode_type, 16#05#),
      1903 => to_slv(opcode_type, 16#0A#),
      1904 => to_slv(opcode_type, 16#10#),
      1905 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#09#),
      1921 => to_slv(opcode_type, 16#09#),
      1922 => to_slv(opcode_type, 16#01#),
      1923 => to_slv(opcode_type, 16#03#),
      1924 => to_slv(opcode_type, 16#11#),
      1925 => to_slv(opcode_type, 16#07#),
      1926 => to_slv(opcode_type, 16#02#),
      1927 => to_slv(opcode_type, 16#10#),
      1928 => to_slv(opcode_type, 16#04#),
      1929 => to_slv(opcode_type, 16#0D#),
      1930 => to_slv(opcode_type, 16#05#),
      1931 => to_slv(opcode_type, 16#07#),
      1932 => to_slv(opcode_type, 16#04#),
      1933 => to_slv(opcode_type, 16#0D#),
      1934 => to_slv(opcode_type, 16#08#),
      1935 => to_slv(opcode_type, 16#0C#),
      1936 => to_slv(opcode_type, 16#11#),
      1937 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#07#),
      1953 => to_slv(opcode_type, 16#07#),
      1954 => to_slv(opcode_type, 16#01#),
      1955 => to_slv(opcode_type, 16#05#),
      1956 => to_slv(opcode_type, 16#0A#),
      1957 => to_slv(opcode_type, 16#08#),
      1958 => to_slv(opcode_type, 16#07#),
      1959 => to_slv(opcode_type, 16#11#),
      1960 => to_slv(opcode_type, 16#0A#),
      1961 => to_slv(opcode_type, 16#03#),
      1962 => to_slv(opcode_type, 16#0C#),
      1963 => to_slv(opcode_type, 16#02#),
      1964 => to_slv(opcode_type, 16#09#),
      1965 => to_slv(opcode_type, 16#07#),
      1966 => to_slv(opcode_type, 16#9E#),
      1967 => to_slv(opcode_type, 16#20#),
      1968 => to_slv(opcode_type, 16#0F#),
      1969 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#06#),
      1985 => to_slv(opcode_type, 16#01#),
      1986 => to_slv(opcode_type, 16#07#),
      1987 => to_slv(opcode_type, 16#04#),
      1988 => to_slv(opcode_type, 16#0F#),
      1989 => to_slv(opcode_type, 16#06#),
      1990 => to_slv(opcode_type, 16#10#),
      1991 => to_slv(opcode_type, 16#0A#),
      1992 => to_slv(opcode_type, 16#07#),
      1993 => to_slv(opcode_type, 16#08#),
      1994 => to_slv(opcode_type, 16#06#),
      1995 => to_slv(opcode_type, 16#10#),
      1996 => to_slv(opcode_type, 16#10#),
      1997 => to_slv(opcode_type, 16#06#),
      1998 => to_slv(opcode_type, 16#0E#),
      1999 => to_slv(opcode_type, 16#0A#),
      2000 => to_slv(opcode_type, 16#E6#),
      2001 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#09#),
      2017 => to_slv(opcode_type, 16#01#),
      2018 => to_slv(opcode_type, 16#03#),
      2019 => to_slv(opcode_type, 16#02#),
      2020 => to_slv(opcode_type, 16#0D#),
      2021 => to_slv(opcode_type, 16#06#),
      2022 => to_slv(opcode_type, 16#06#),
      2023 => to_slv(opcode_type, 16#03#),
      2024 => to_slv(opcode_type, 16#0C#),
      2025 => to_slv(opcode_type, 16#02#),
      2026 => to_slv(opcode_type, 16#0A#),
      2027 => to_slv(opcode_type, 16#06#),
      2028 => to_slv(opcode_type, 16#08#),
      2029 => to_slv(opcode_type, 16#AF#),
      2030 => to_slv(opcode_type, 16#60#),
      2031 => to_slv(opcode_type, 16#05#),
      2032 => to_slv(opcode_type, 16#11#),
      2033 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#07#),
      2049 => to_slv(opcode_type, 16#08#),
      2050 => to_slv(opcode_type, 16#04#),
      2051 => to_slv(opcode_type, 16#03#),
      2052 => to_slv(opcode_type, 16#0B#),
      2053 => to_slv(opcode_type, 16#01#),
      2054 => to_slv(opcode_type, 16#02#),
      2055 => to_slv(opcode_type, 16#0E#),
      2056 => to_slv(opcode_type, 16#08#),
      2057 => to_slv(opcode_type, 16#04#),
      2058 => to_slv(opcode_type, 16#08#),
      2059 => to_slv(opcode_type, 16#0E#),
      2060 => to_slv(opcode_type, 16#10#),
      2061 => to_slv(opcode_type, 16#05#),
      2062 => to_slv(opcode_type, 16#06#),
      2063 => to_slv(opcode_type, 16#0C#),
      2064 => to_slv(opcode_type, 16#10#),
      2065 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#08#),
      2081 => to_slv(opcode_type, 16#07#),
      2082 => to_slv(opcode_type, 16#06#),
      2083 => to_slv(opcode_type, 16#02#),
      2084 => to_slv(opcode_type, 16#0A#),
      2085 => to_slv(opcode_type, 16#02#),
      2086 => to_slv(opcode_type, 16#11#),
      2087 => to_slv(opcode_type, 16#04#),
      2088 => to_slv(opcode_type, 16#03#),
      2089 => to_slv(opcode_type, 16#0B#),
      2090 => to_slv(opcode_type, 16#03#),
      2091 => to_slv(opcode_type, 16#07#),
      2092 => to_slv(opcode_type, 16#06#),
      2093 => to_slv(opcode_type, 16#0E#),
      2094 => to_slv(opcode_type, 16#0D#),
      2095 => to_slv(opcode_type, 16#03#),
      2096 => to_slv(opcode_type, 16#0B#),
      2097 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#06#),
      2113 => to_slv(opcode_type, 16#09#),
      2114 => to_slv(opcode_type, 16#03#),
      2115 => to_slv(opcode_type, 16#05#),
      2116 => to_slv(opcode_type, 16#10#),
      2117 => to_slv(opcode_type, 16#03#),
      2118 => to_slv(opcode_type, 16#05#),
      2119 => to_slv(opcode_type, 16#0F#),
      2120 => to_slv(opcode_type, 16#07#),
      2121 => to_slv(opcode_type, 16#01#),
      2122 => to_slv(opcode_type, 16#05#),
      2123 => to_slv(opcode_type, 16#0D#),
      2124 => to_slv(opcode_type, 16#06#),
      2125 => to_slv(opcode_type, 16#01#),
      2126 => to_slv(opcode_type, 16#11#),
      2127 => to_slv(opcode_type, 16#03#),
      2128 => to_slv(opcode_type, 16#0B#),
      2129 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#07#),
      2145 => to_slv(opcode_type, 16#01#),
      2146 => to_slv(opcode_type, 16#08#),
      2147 => to_slv(opcode_type, 16#08#),
      2148 => to_slv(opcode_type, 16#11#),
      2149 => to_slv(opcode_type, 16#0C#),
      2150 => to_slv(opcode_type, 16#03#),
      2151 => to_slv(opcode_type, 16#0F#),
      2152 => to_slv(opcode_type, 16#06#),
      2153 => to_slv(opcode_type, 16#03#),
      2154 => to_slv(opcode_type, 16#09#),
      2155 => to_slv(opcode_type, 16#0C#),
      2156 => to_slv(opcode_type, 16#10#),
      2157 => to_slv(opcode_type, 16#02#),
      2158 => to_slv(opcode_type, 16#07#),
      2159 => to_slv(opcode_type, 16#11#),
      2160 => to_slv(opcode_type, 16#0E#),
      2161 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#09#),
      2177 => to_slv(opcode_type, 16#03#),
      2178 => to_slv(opcode_type, 16#06#),
      2179 => to_slv(opcode_type, 16#05#),
      2180 => to_slv(opcode_type, 16#0E#),
      2181 => to_slv(opcode_type, 16#05#),
      2182 => to_slv(opcode_type, 16#0F#),
      2183 => to_slv(opcode_type, 16#09#),
      2184 => to_slv(opcode_type, 16#03#),
      2185 => to_slv(opcode_type, 16#08#),
      2186 => to_slv(opcode_type, 16#10#),
      2187 => to_slv(opcode_type, 16#E7#),
      2188 => to_slv(opcode_type, 16#07#),
      2189 => to_slv(opcode_type, 16#06#),
      2190 => to_slv(opcode_type, 16#0D#),
      2191 => to_slv(opcode_type, 16#AD#),
      2192 => to_slv(opcode_type, 16#0A#),
      2193 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#06#),
      2209 => to_slv(opcode_type, 16#04#),
      2210 => to_slv(opcode_type, 16#05#),
      2211 => to_slv(opcode_type, 16#07#),
      2212 => to_slv(opcode_type, 16#10#),
      2213 => to_slv(opcode_type, 16#10#),
      2214 => to_slv(opcode_type, 16#06#),
      2215 => to_slv(opcode_type, 16#02#),
      2216 => to_slv(opcode_type, 16#02#),
      2217 => to_slv(opcode_type, 16#11#),
      2218 => to_slv(opcode_type, 16#07#),
      2219 => to_slv(opcode_type, 16#09#),
      2220 => to_slv(opcode_type, 16#0C#),
      2221 => to_slv(opcode_type, 16#0C#),
      2222 => to_slv(opcode_type, 16#08#),
      2223 => to_slv(opcode_type, 16#0C#),
      2224 => to_slv(opcode_type, 16#0D#),
      2225 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#08#),
      2241 => to_slv(opcode_type, 16#01#),
      2242 => to_slv(opcode_type, 16#04#),
      2243 => to_slv(opcode_type, 16#04#),
      2244 => to_slv(opcode_type, 16#0C#),
      2245 => to_slv(opcode_type, 16#09#),
      2246 => to_slv(opcode_type, 16#03#),
      2247 => to_slv(opcode_type, 16#06#),
      2248 => to_slv(opcode_type, 16#A5#),
      2249 => to_slv(opcode_type, 16#0E#),
      2250 => to_slv(opcode_type, 16#09#),
      2251 => to_slv(opcode_type, 16#09#),
      2252 => to_slv(opcode_type, 16#0F#),
      2253 => to_slv(opcode_type, 16#5D#),
      2254 => to_slv(opcode_type, 16#06#),
      2255 => to_slv(opcode_type, 16#0B#),
      2256 => to_slv(opcode_type, 16#0F#),
      2257 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#09#),
      2273 => to_slv(opcode_type, 16#09#),
      2274 => to_slv(opcode_type, 16#09#),
      2275 => to_slv(opcode_type, 16#01#),
      2276 => to_slv(opcode_type, 16#11#),
      2277 => to_slv(opcode_type, 16#02#),
      2278 => to_slv(opcode_type, 16#11#),
      2279 => to_slv(opcode_type, 16#07#),
      2280 => to_slv(opcode_type, 16#08#),
      2281 => to_slv(opcode_type, 16#10#),
      2282 => to_slv(opcode_type, 16#31#),
      2283 => to_slv(opcode_type, 16#03#),
      2284 => to_slv(opcode_type, 16#0A#),
      2285 => to_slv(opcode_type, 16#02#),
      2286 => to_slv(opcode_type, 16#04#),
      2287 => to_slv(opcode_type, 16#04#),
      2288 => to_slv(opcode_type, 16#11#),
      2289 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#07#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#06#),
      2307 => to_slv(opcode_type, 16#01#),
      2308 => to_slv(opcode_type, 16#D8#),
      2309 => to_slv(opcode_type, 16#07#),
      2310 => to_slv(opcode_type, 16#0C#),
      2311 => to_slv(opcode_type, 16#0C#),
      2312 => to_slv(opcode_type, 16#05#),
      2313 => to_slv(opcode_type, 16#08#),
      2314 => to_slv(opcode_type, 16#0C#),
      2315 => to_slv(opcode_type, 16#0D#),
      2316 => to_slv(opcode_type, 16#09#),
      2317 => to_slv(opcode_type, 16#01#),
      2318 => to_slv(opcode_type, 16#03#),
      2319 => to_slv(opcode_type, 16#0B#),
      2320 => to_slv(opcode_type, 16#10#),
      2321 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#08#),
      2337 => to_slv(opcode_type, 16#03#),
      2338 => to_slv(opcode_type, 16#03#),
      2339 => to_slv(opcode_type, 16#04#),
      2340 => to_slv(opcode_type, 16#0C#),
      2341 => to_slv(opcode_type, 16#06#),
      2342 => to_slv(opcode_type, 16#02#),
      2343 => to_slv(opcode_type, 16#08#),
      2344 => to_slv(opcode_type, 16#11#),
      2345 => to_slv(opcode_type, 16#0C#),
      2346 => to_slv(opcode_type, 16#09#),
      2347 => to_slv(opcode_type, 16#07#),
      2348 => to_slv(opcode_type, 16#0D#),
      2349 => to_slv(opcode_type, 16#0B#),
      2350 => to_slv(opcode_type, 16#06#),
      2351 => to_slv(opcode_type, 16#0D#),
      2352 => to_slv(opcode_type, 16#0F#),
      2353 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#07#),
      2369 => to_slv(opcode_type, 16#03#),
      2370 => to_slv(opcode_type, 16#05#),
      2371 => to_slv(opcode_type, 16#01#),
      2372 => to_slv(opcode_type, 16#0A#),
      2373 => to_slv(opcode_type, 16#07#),
      2374 => to_slv(opcode_type, 16#09#),
      2375 => to_slv(opcode_type, 16#02#),
      2376 => to_slv(opcode_type, 16#0B#),
      2377 => to_slv(opcode_type, 16#04#),
      2378 => to_slv(opcode_type, 16#0E#),
      2379 => to_slv(opcode_type, 16#06#),
      2380 => to_slv(opcode_type, 16#03#),
      2381 => to_slv(opcode_type, 16#0D#),
      2382 => to_slv(opcode_type, 16#06#),
      2383 => to_slv(opcode_type, 16#0E#),
      2384 => to_slv(opcode_type, 16#0D#),
      2385 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#08#),
      2401 => to_slv(opcode_type, 16#07#),
      2402 => to_slv(opcode_type, 16#02#),
      2403 => to_slv(opcode_type, 16#04#),
      2404 => to_slv(opcode_type, 16#11#),
      2405 => to_slv(opcode_type, 16#03#),
      2406 => to_slv(opcode_type, 16#02#),
      2407 => to_slv(opcode_type, 16#0D#),
      2408 => to_slv(opcode_type, 16#06#),
      2409 => to_slv(opcode_type, 16#04#),
      2410 => to_slv(opcode_type, 16#07#),
      2411 => to_slv(opcode_type, 16#0A#),
      2412 => to_slv(opcode_type, 16#F1#),
      2413 => to_slv(opcode_type, 16#08#),
      2414 => to_slv(opcode_type, 16#03#),
      2415 => to_slv(opcode_type, 16#10#),
      2416 => to_slv(opcode_type, 16#0E#),
      2417 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#08#),
      2433 => to_slv(opcode_type, 16#03#),
      2434 => to_slv(opcode_type, 16#09#),
      2435 => to_slv(opcode_type, 16#03#),
      2436 => to_slv(opcode_type, 16#0B#),
      2437 => to_slv(opcode_type, 16#04#),
      2438 => to_slv(opcode_type, 16#0C#),
      2439 => to_slv(opcode_type, 16#06#),
      2440 => to_slv(opcode_type, 16#03#),
      2441 => to_slv(opcode_type, 16#07#),
      2442 => to_slv(opcode_type, 16#0C#),
      2443 => to_slv(opcode_type, 16#0A#),
      2444 => to_slv(opcode_type, 16#07#),
      2445 => to_slv(opcode_type, 16#02#),
      2446 => to_slv(opcode_type, 16#11#),
      2447 => to_slv(opcode_type, 16#01#),
      2448 => to_slv(opcode_type, 16#0A#),
      2449 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#06#),
      2465 => to_slv(opcode_type, 16#02#),
      2466 => to_slv(opcode_type, 16#06#),
      2467 => to_slv(opcode_type, 16#01#),
      2468 => to_slv(opcode_type, 16#0C#),
      2469 => to_slv(opcode_type, 16#08#),
      2470 => to_slv(opcode_type, 16#85#),
      2471 => to_slv(opcode_type, 16#0F#),
      2472 => to_slv(opcode_type, 16#07#),
      2473 => to_slv(opcode_type, 16#01#),
      2474 => to_slv(opcode_type, 16#07#),
      2475 => to_slv(opcode_type, 16#F8#),
      2476 => to_slv(opcode_type, 16#0A#),
      2477 => to_slv(opcode_type, 16#03#),
      2478 => to_slv(opcode_type, 16#08#),
      2479 => to_slv(opcode_type, 16#0D#),
      2480 => to_slv(opcode_type, 16#0B#),
      2481 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#06#),
      2497 => to_slv(opcode_type, 16#03#),
      2498 => to_slv(opcode_type, 16#02#),
      2499 => to_slv(opcode_type, 16#02#),
      2500 => to_slv(opcode_type, 16#6B#),
      2501 => to_slv(opcode_type, 16#09#),
      2502 => to_slv(opcode_type, 16#06#),
      2503 => to_slv(opcode_type, 16#09#),
      2504 => to_slv(opcode_type, 16#11#),
      2505 => to_slv(opcode_type, 16#11#),
      2506 => to_slv(opcode_type, 16#07#),
      2507 => to_slv(opcode_type, 16#0A#),
      2508 => to_slv(opcode_type, 16#0D#),
      2509 => to_slv(opcode_type, 16#02#),
      2510 => to_slv(opcode_type, 16#09#),
      2511 => to_slv(opcode_type, 16#50#),
      2512 => to_slv(opcode_type, 16#0A#),
      2513 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#04#),
      2530 => to_slv(opcode_type, 16#08#),
      2531 => to_slv(opcode_type, 16#03#),
      2532 => to_slv(opcode_type, 16#11#),
      2533 => to_slv(opcode_type, 16#02#),
      2534 => to_slv(opcode_type, 16#0F#),
      2535 => to_slv(opcode_type, 16#07#),
      2536 => to_slv(opcode_type, 16#09#),
      2537 => to_slv(opcode_type, 16#01#),
      2538 => to_slv(opcode_type, 16#0C#),
      2539 => to_slv(opcode_type, 16#07#),
      2540 => to_slv(opcode_type, 16#0F#),
      2541 => to_slv(opcode_type, 16#11#),
      2542 => to_slv(opcode_type, 16#03#),
      2543 => to_slv(opcode_type, 16#02#),
      2544 => to_slv(opcode_type, 16#0D#),
      2545 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#08#),
      2561 => to_slv(opcode_type, 16#03#),
      2562 => to_slv(opcode_type, 16#01#),
      2563 => to_slv(opcode_type, 16#06#),
      2564 => to_slv(opcode_type, 16#76#),
      2565 => to_slv(opcode_type, 16#AA#),
      2566 => to_slv(opcode_type, 16#09#),
      2567 => to_slv(opcode_type, 16#03#),
      2568 => to_slv(opcode_type, 16#05#),
      2569 => to_slv(opcode_type, 16#0E#),
      2570 => to_slv(opcode_type, 16#06#),
      2571 => to_slv(opcode_type, 16#09#),
      2572 => to_slv(opcode_type, 16#0A#),
      2573 => to_slv(opcode_type, 16#10#),
      2574 => to_slv(opcode_type, 16#06#),
      2575 => to_slv(opcode_type, 16#0F#),
      2576 => to_slv(opcode_type, 16#0E#),
      2577 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#09#),
      2593 => to_slv(opcode_type, 16#08#),
      2594 => to_slv(opcode_type, 16#03#),
      2595 => to_slv(opcode_type, 16#08#),
      2596 => to_slv(opcode_type, 16#0E#),
      2597 => to_slv(opcode_type, 16#0D#),
      2598 => to_slv(opcode_type, 16#05#),
      2599 => to_slv(opcode_type, 16#01#),
      2600 => to_slv(opcode_type, 16#0F#),
      2601 => to_slv(opcode_type, 16#08#),
      2602 => to_slv(opcode_type, 16#09#),
      2603 => to_slv(opcode_type, 16#03#),
      2604 => to_slv(opcode_type, 16#0B#),
      2605 => to_slv(opcode_type, 16#04#),
      2606 => to_slv(opcode_type, 16#0B#),
      2607 => to_slv(opcode_type, 16#02#),
      2608 => to_slv(opcode_type, 16#11#),
      2609 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#06#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#07#),
      2627 => to_slv(opcode_type, 16#04#),
      2628 => to_slv(opcode_type, 16#10#),
      2629 => to_slv(opcode_type, 16#08#),
      2630 => to_slv(opcode_type, 16#0B#),
      2631 => to_slv(opcode_type, 16#A5#),
      2632 => to_slv(opcode_type, 16#08#),
      2633 => to_slv(opcode_type, 16#02#),
      2634 => to_slv(opcode_type, 16#10#),
      2635 => to_slv(opcode_type, 16#08#),
      2636 => to_slv(opcode_type, 16#11#),
      2637 => to_slv(opcode_type, 16#0A#),
      2638 => to_slv(opcode_type, 16#01#),
      2639 => to_slv(opcode_type, 16#04#),
      2640 => to_slv(opcode_type, 16#0A#),
      2641 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#08#),
      2657 => to_slv(opcode_type, 16#09#),
      2658 => to_slv(opcode_type, 16#07#),
      2659 => to_slv(opcode_type, 16#02#),
      2660 => to_slv(opcode_type, 16#FE#),
      2661 => to_slv(opcode_type, 16#03#),
      2662 => to_slv(opcode_type, 16#9F#),
      2663 => to_slv(opcode_type, 16#08#),
      2664 => to_slv(opcode_type, 16#06#),
      2665 => to_slv(opcode_type, 16#EF#),
      2666 => to_slv(opcode_type, 16#0F#),
      2667 => to_slv(opcode_type, 16#05#),
      2668 => to_slv(opcode_type, 16#11#),
      2669 => to_slv(opcode_type, 16#07#),
      2670 => to_slv(opcode_type, 16#02#),
      2671 => to_slv(opcode_type, 16#0F#),
      2672 => to_slv(opcode_type, 16#0F#),
      2673 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#06#),
      2689 => to_slv(opcode_type, 16#07#),
      2690 => to_slv(opcode_type, 16#02#),
      2691 => to_slv(opcode_type, 16#03#),
      2692 => to_slv(opcode_type, 16#0A#),
      2693 => to_slv(opcode_type, 16#05#),
      2694 => to_slv(opcode_type, 16#08#),
      2695 => to_slv(opcode_type, 16#0D#),
      2696 => to_slv(opcode_type, 16#0E#),
      2697 => to_slv(opcode_type, 16#02#),
      2698 => to_slv(opcode_type, 16#06#),
      2699 => to_slv(opcode_type, 16#08#),
      2700 => to_slv(opcode_type, 16#0A#),
      2701 => to_slv(opcode_type, 16#0F#),
      2702 => to_slv(opcode_type, 16#07#),
      2703 => to_slv(opcode_type, 16#0B#),
      2704 => to_slv(opcode_type, 16#10#),
      2705 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#06#),
      2721 => to_slv(opcode_type, 16#02#),
      2722 => to_slv(opcode_type, 16#02#),
      2723 => to_slv(opcode_type, 16#09#),
      2724 => to_slv(opcode_type, 16#10#),
      2725 => to_slv(opcode_type, 16#0D#),
      2726 => to_slv(opcode_type, 16#06#),
      2727 => to_slv(opcode_type, 16#07#),
      2728 => to_slv(opcode_type, 16#03#),
      2729 => to_slv(opcode_type, 16#0F#),
      2730 => to_slv(opcode_type, 16#03#),
      2731 => to_slv(opcode_type, 16#0A#),
      2732 => to_slv(opcode_type, 16#07#),
      2733 => to_slv(opcode_type, 16#07#),
      2734 => to_slv(opcode_type, 16#0F#),
      2735 => to_slv(opcode_type, 16#0B#),
      2736 => to_slv(opcode_type, 16#10#),
      2737 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#06#),
      2753 => to_slv(opcode_type, 16#03#),
      2754 => to_slv(opcode_type, 16#05#),
      2755 => to_slv(opcode_type, 16#07#),
      2756 => to_slv(opcode_type, 16#11#),
      2757 => to_slv(opcode_type, 16#10#),
      2758 => to_slv(opcode_type, 16#07#),
      2759 => to_slv(opcode_type, 16#01#),
      2760 => to_slv(opcode_type, 16#08#),
      2761 => to_slv(opcode_type, 16#0F#),
      2762 => to_slv(opcode_type, 16#11#),
      2763 => to_slv(opcode_type, 16#06#),
      2764 => to_slv(opcode_type, 16#04#),
      2765 => to_slv(opcode_type, 16#0A#),
      2766 => to_slv(opcode_type, 16#06#),
      2767 => to_slv(opcode_type, 16#0A#),
      2768 => to_slv(opcode_type, 16#BD#),
      2769 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#07#),
      2785 => to_slv(opcode_type, 16#06#),
      2786 => to_slv(opcode_type, 16#02#),
      2787 => to_slv(opcode_type, 16#08#),
      2788 => to_slv(opcode_type, 16#0F#),
      2789 => to_slv(opcode_type, 16#10#),
      2790 => to_slv(opcode_type, 16#09#),
      2791 => to_slv(opcode_type, 16#04#),
      2792 => to_slv(opcode_type, 16#0F#),
      2793 => to_slv(opcode_type, 16#01#),
      2794 => to_slv(opcode_type, 16#0C#),
      2795 => to_slv(opcode_type, 16#06#),
      2796 => to_slv(opcode_type, 16#05#),
      2797 => to_slv(opcode_type, 16#05#),
      2798 => to_slv(opcode_type, 16#0A#),
      2799 => to_slv(opcode_type, 16#05#),
      2800 => to_slv(opcode_type, 16#11#),
      2801 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#07#),
      2817 => to_slv(opcode_type, 16#08#),
      2818 => to_slv(opcode_type, 16#06#),
      2819 => to_slv(opcode_type, 16#07#),
      2820 => to_slv(opcode_type, 16#0A#),
      2821 => to_slv(opcode_type, 16#0F#),
      2822 => to_slv(opcode_type, 16#01#),
      2823 => to_slv(opcode_type, 16#0F#),
      2824 => to_slv(opcode_type, 16#06#),
      2825 => to_slv(opcode_type, 16#05#),
      2826 => to_slv(opcode_type, 16#10#),
      2827 => to_slv(opcode_type, 16#05#),
      2828 => to_slv(opcode_type, 16#0F#),
      2829 => to_slv(opcode_type, 16#05#),
      2830 => to_slv(opcode_type, 16#08#),
      2831 => to_slv(opcode_type, 16#0E#),
      2832 => to_slv(opcode_type, 16#0F#),
      2833 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#06#),
      2849 => to_slv(opcode_type, 16#08#),
      2850 => to_slv(opcode_type, 16#03#),
      2851 => to_slv(opcode_type, 16#06#),
      2852 => to_slv(opcode_type, 16#0E#),
      2853 => to_slv(opcode_type, 16#0F#),
      2854 => to_slv(opcode_type, 16#05#),
      2855 => to_slv(opcode_type, 16#03#),
      2856 => to_slv(opcode_type, 16#0C#),
      2857 => to_slv(opcode_type, 16#08#),
      2858 => to_slv(opcode_type, 16#08#),
      2859 => to_slv(opcode_type, 16#06#),
      2860 => to_slv(opcode_type, 16#0B#),
      2861 => to_slv(opcode_type, 16#0F#),
      2862 => to_slv(opcode_type, 16#05#),
      2863 => to_slv(opcode_type, 16#0B#),
      2864 => to_slv(opcode_type, 16#0A#),
      2865 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#09#),
      2881 => to_slv(opcode_type, 16#04#),
      2882 => to_slv(opcode_type, 16#08#),
      2883 => to_slv(opcode_type, 16#05#),
      2884 => to_slv(opcode_type, 16#0A#),
      2885 => to_slv(opcode_type, 16#06#),
      2886 => to_slv(opcode_type, 16#0E#),
      2887 => to_slv(opcode_type, 16#0F#),
      2888 => to_slv(opcode_type, 16#06#),
      2889 => to_slv(opcode_type, 16#05#),
      2890 => to_slv(opcode_type, 16#07#),
      2891 => to_slv(opcode_type, 16#0E#),
      2892 => to_slv(opcode_type, 16#0B#),
      2893 => to_slv(opcode_type, 16#05#),
      2894 => to_slv(opcode_type, 16#07#),
      2895 => to_slv(opcode_type, 16#0F#),
      2896 => to_slv(opcode_type, 16#10#),
      2897 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#06#),
      2913 => to_slv(opcode_type, 16#03#),
      2914 => to_slv(opcode_type, 16#06#),
      2915 => to_slv(opcode_type, 16#05#),
      2916 => to_slv(opcode_type, 16#0D#),
      2917 => to_slv(opcode_type, 16#04#),
      2918 => to_slv(opcode_type, 16#D3#),
      2919 => to_slv(opcode_type, 16#07#),
      2920 => to_slv(opcode_type, 16#06#),
      2921 => to_slv(opcode_type, 16#04#),
      2922 => to_slv(opcode_type, 16#CE#),
      2923 => to_slv(opcode_type, 16#07#),
      2924 => to_slv(opcode_type, 16#0A#),
      2925 => to_slv(opcode_type, 16#0E#),
      2926 => to_slv(opcode_type, 16#08#),
      2927 => to_slv(opcode_type, 16#0E#),
      2928 => to_slv(opcode_type, 16#11#),
      2929 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#08#),
      2945 => to_slv(opcode_type, 16#09#),
      2946 => to_slv(opcode_type, 16#05#),
      2947 => to_slv(opcode_type, 16#09#),
      2948 => to_slv(opcode_type, 16#0C#),
      2949 => to_slv(opcode_type, 16#0A#),
      2950 => to_slv(opcode_type, 16#07#),
      2951 => to_slv(opcode_type, 16#03#),
      2952 => to_slv(opcode_type, 16#C2#),
      2953 => to_slv(opcode_type, 16#02#),
      2954 => to_slv(opcode_type, 16#0F#),
      2955 => to_slv(opcode_type, 16#01#),
      2956 => to_slv(opcode_type, 16#09#),
      2957 => to_slv(opcode_type, 16#03#),
      2958 => to_slv(opcode_type, 16#0F#),
      2959 => to_slv(opcode_type, 16#03#),
      2960 => to_slv(opcode_type, 16#C8#),
      2961 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#07#),
      2977 => to_slv(opcode_type, 16#03#),
      2978 => to_slv(opcode_type, 16#08#),
      2979 => to_slv(opcode_type, 16#04#),
      2980 => to_slv(opcode_type, 16#0B#),
      2981 => to_slv(opcode_type, 16#04#),
      2982 => to_slv(opcode_type, 16#0C#),
      2983 => to_slv(opcode_type, 16#06#),
      2984 => to_slv(opcode_type, 16#09#),
      2985 => to_slv(opcode_type, 16#01#),
      2986 => to_slv(opcode_type, 16#0C#),
      2987 => to_slv(opcode_type, 16#07#),
      2988 => to_slv(opcode_type, 16#11#),
      2989 => to_slv(opcode_type, 16#5F#),
      2990 => to_slv(opcode_type, 16#04#),
      2991 => to_slv(opcode_type, 16#03#),
      2992 => to_slv(opcode_type, 16#11#),
      2993 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#07#),
      3009 => to_slv(opcode_type, 16#04#),
      3010 => to_slv(opcode_type, 16#06#),
      3011 => to_slv(opcode_type, 16#06#),
      3012 => to_slv(opcode_type, 16#62#),
      3013 => to_slv(opcode_type, 16#72#),
      3014 => to_slv(opcode_type, 16#08#),
      3015 => to_slv(opcode_type, 16#0B#),
      3016 => to_slv(opcode_type, 16#0C#),
      3017 => to_slv(opcode_type, 16#09#),
      3018 => to_slv(opcode_type, 16#08#),
      3019 => to_slv(opcode_type, 16#02#),
      3020 => to_slv(opcode_type, 16#11#),
      3021 => to_slv(opcode_type, 16#02#),
      3022 => to_slv(opcode_type, 16#0C#),
      3023 => to_slv(opcode_type, 16#05#),
      3024 => to_slv(opcode_type, 16#0A#),
      3025 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#07#),
      3041 => to_slv(opcode_type, 16#09#),
      3042 => to_slv(opcode_type, 16#04#),
      3043 => to_slv(opcode_type, 16#04#),
      3044 => to_slv(opcode_type, 16#10#),
      3045 => to_slv(opcode_type, 16#04#),
      3046 => to_slv(opcode_type, 16#02#),
      3047 => to_slv(opcode_type, 16#0F#),
      3048 => to_slv(opcode_type, 16#06#),
      3049 => to_slv(opcode_type, 16#01#),
      3050 => to_slv(opcode_type, 16#03#),
      3051 => to_slv(opcode_type, 16#11#),
      3052 => to_slv(opcode_type, 16#06#),
      3053 => to_slv(opcode_type, 16#03#),
      3054 => to_slv(opcode_type, 16#1B#),
      3055 => to_slv(opcode_type, 16#02#),
      3056 => to_slv(opcode_type, 16#10#),
      3057 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#08#),
      3073 => to_slv(opcode_type, 16#08#),
      3074 => to_slv(opcode_type, 16#09#),
      3075 => to_slv(opcode_type, 16#09#),
      3076 => to_slv(opcode_type, 16#0F#),
      3077 => to_slv(opcode_type, 16#E0#),
      3078 => to_slv(opcode_type, 16#01#),
      3079 => to_slv(opcode_type, 16#0D#),
      3080 => to_slv(opcode_type, 16#06#),
      3081 => to_slv(opcode_type, 16#09#),
      3082 => to_slv(opcode_type, 16#0C#),
      3083 => to_slv(opcode_type, 16#0A#),
      3084 => to_slv(opcode_type, 16#09#),
      3085 => to_slv(opcode_type, 16#11#),
      3086 => to_slv(opcode_type, 16#10#),
      3087 => to_slv(opcode_type, 16#03#),
      3088 => to_slv(opcode_type, 16#11#),
      3089 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#09#),
      3105 => to_slv(opcode_type, 16#08#),
      3106 => to_slv(opcode_type, 16#01#),
      3107 => to_slv(opcode_type, 16#09#),
      3108 => to_slv(opcode_type, 16#0A#),
      3109 => to_slv(opcode_type, 16#0C#),
      3110 => to_slv(opcode_type, 16#01#),
      3111 => to_slv(opcode_type, 16#02#),
      3112 => to_slv(opcode_type, 16#0C#),
      3113 => to_slv(opcode_type, 16#01#),
      3114 => to_slv(opcode_type, 16#08#),
      3115 => to_slv(opcode_type, 16#08#),
      3116 => to_slv(opcode_type, 16#0E#),
      3117 => to_slv(opcode_type, 16#0A#),
      3118 => to_slv(opcode_type, 16#06#),
      3119 => to_slv(opcode_type, 16#0B#),
      3120 => to_slv(opcode_type, 16#0A#),
      3121 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#09#),
      3137 => to_slv(opcode_type, 16#05#),
      3138 => to_slv(opcode_type, 16#05#),
      3139 => to_slv(opcode_type, 16#01#),
      3140 => to_slv(opcode_type, 16#0D#),
      3141 => to_slv(opcode_type, 16#06#),
      3142 => to_slv(opcode_type, 16#08#),
      3143 => to_slv(opcode_type, 16#06#),
      3144 => to_slv(opcode_type, 16#0F#),
      3145 => to_slv(opcode_type, 16#0F#),
      3146 => to_slv(opcode_type, 16#05#),
      3147 => to_slv(opcode_type, 16#0B#),
      3148 => to_slv(opcode_type, 16#06#),
      3149 => to_slv(opcode_type, 16#05#),
      3150 => to_slv(opcode_type, 16#0B#),
      3151 => to_slv(opcode_type, 16#03#),
      3152 => to_slv(opcode_type, 16#2C#),
      3153 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#07#),
      3169 => to_slv(opcode_type, 16#08#),
      3170 => to_slv(opcode_type, 16#03#),
      3171 => to_slv(opcode_type, 16#04#),
      3172 => to_slv(opcode_type, 16#0C#),
      3173 => to_slv(opcode_type, 16#09#),
      3174 => to_slv(opcode_type, 16#09#),
      3175 => to_slv(opcode_type, 16#0B#),
      3176 => to_slv(opcode_type, 16#0F#),
      3177 => to_slv(opcode_type, 16#09#),
      3178 => to_slv(opcode_type, 16#10#),
      3179 => to_slv(opcode_type, 16#0C#),
      3180 => to_slv(opcode_type, 16#02#),
      3181 => to_slv(opcode_type, 16#05#),
      3182 => to_slv(opcode_type, 16#06#),
      3183 => to_slv(opcode_type, 16#0D#),
      3184 => to_slv(opcode_type, 16#0D#),
      3185 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#06#),
      3201 => to_slv(opcode_type, 16#04#),
      3202 => to_slv(opcode_type, 16#02#),
      3203 => to_slv(opcode_type, 16#05#),
      3204 => to_slv(opcode_type, 16#11#),
      3205 => to_slv(opcode_type, 16#06#),
      3206 => to_slv(opcode_type, 16#05#),
      3207 => to_slv(opcode_type, 16#07#),
      3208 => to_slv(opcode_type, 16#0E#),
      3209 => to_slv(opcode_type, 16#0D#),
      3210 => to_slv(opcode_type, 16#06#),
      3211 => to_slv(opcode_type, 16#06#),
      3212 => to_slv(opcode_type, 16#0B#),
      3213 => to_slv(opcode_type, 16#11#),
      3214 => to_slv(opcode_type, 16#08#),
      3215 => to_slv(opcode_type, 16#10#),
      3216 => to_slv(opcode_type, 16#0B#),
      3217 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#02#),
      3234 => to_slv(opcode_type, 16#08#),
      3235 => to_slv(opcode_type, 16#01#),
      3236 => to_slv(opcode_type, 16#0F#),
      3237 => to_slv(opcode_type, 16#02#),
      3238 => to_slv(opcode_type, 16#1C#),
      3239 => to_slv(opcode_type, 16#09#),
      3240 => to_slv(opcode_type, 16#07#),
      3241 => to_slv(opcode_type, 16#05#),
      3242 => to_slv(opcode_type, 16#0F#),
      3243 => to_slv(opcode_type, 16#08#),
      3244 => to_slv(opcode_type, 16#10#),
      3245 => to_slv(opcode_type, 16#0E#),
      3246 => to_slv(opcode_type, 16#05#),
      3247 => to_slv(opcode_type, 16#01#),
      3248 => to_slv(opcode_type, 16#11#),
      3249 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#08#),
      3265 => to_slv(opcode_type, 16#05#),
      3266 => to_slv(opcode_type, 16#05#),
      3267 => to_slv(opcode_type, 16#08#),
      3268 => to_slv(opcode_type, 16#0E#),
      3269 => to_slv(opcode_type, 16#0A#),
      3270 => to_slv(opcode_type, 16#08#),
      3271 => to_slv(opcode_type, 16#04#),
      3272 => to_slv(opcode_type, 16#06#),
      3273 => to_slv(opcode_type, 16#0C#),
      3274 => to_slv(opcode_type, 16#6F#),
      3275 => to_slv(opcode_type, 16#07#),
      3276 => to_slv(opcode_type, 16#09#),
      3277 => to_slv(opcode_type, 16#0D#),
      3278 => to_slv(opcode_type, 16#11#),
      3279 => to_slv(opcode_type, 16#05#),
      3280 => to_slv(opcode_type, 16#0D#),
      3281 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#09#),
      3297 => to_slv(opcode_type, 16#02#),
      3298 => to_slv(opcode_type, 16#08#),
      3299 => to_slv(opcode_type, 16#01#),
      3300 => to_slv(opcode_type, 16#0B#),
      3301 => to_slv(opcode_type, 16#03#),
      3302 => to_slv(opcode_type, 16#0F#),
      3303 => to_slv(opcode_type, 16#08#),
      3304 => to_slv(opcode_type, 16#09#),
      3305 => to_slv(opcode_type, 16#08#),
      3306 => to_slv(opcode_type, 16#0A#),
      3307 => to_slv(opcode_type, 16#0B#),
      3308 => to_slv(opcode_type, 16#06#),
      3309 => to_slv(opcode_type, 16#0D#),
      3310 => to_slv(opcode_type, 16#0B#),
      3311 => to_slv(opcode_type, 16#01#),
      3312 => to_slv(opcode_type, 16#0A#),
      3313 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#08#),
      3329 => to_slv(opcode_type, 16#01#),
      3330 => to_slv(opcode_type, 16#03#),
      3331 => to_slv(opcode_type, 16#03#),
      3332 => to_slv(opcode_type, 16#0B#),
      3333 => to_slv(opcode_type, 16#08#),
      3334 => to_slv(opcode_type, 16#05#),
      3335 => to_slv(opcode_type, 16#06#),
      3336 => to_slv(opcode_type, 16#0A#),
      3337 => to_slv(opcode_type, 16#10#),
      3338 => to_slv(opcode_type, 16#07#),
      3339 => to_slv(opcode_type, 16#08#),
      3340 => to_slv(opcode_type, 16#0A#),
      3341 => to_slv(opcode_type, 16#0B#),
      3342 => to_slv(opcode_type, 16#07#),
      3343 => to_slv(opcode_type, 16#11#),
      3344 => to_slv(opcode_type, 16#0D#),
      3345 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#06#),
      3361 => to_slv(opcode_type, 16#03#),
      3362 => to_slv(opcode_type, 16#06#),
      3363 => to_slv(opcode_type, 16#05#),
      3364 => to_slv(opcode_type, 16#0A#),
      3365 => to_slv(opcode_type, 16#04#),
      3366 => to_slv(opcode_type, 16#0B#),
      3367 => to_slv(opcode_type, 16#09#),
      3368 => to_slv(opcode_type, 16#05#),
      3369 => to_slv(opcode_type, 16#06#),
      3370 => to_slv(opcode_type, 16#0D#),
      3371 => to_slv(opcode_type, 16#0F#),
      3372 => to_slv(opcode_type, 16#06#),
      3373 => to_slv(opcode_type, 16#08#),
      3374 => to_slv(opcode_type, 16#0F#),
      3375 => to_slv(opcode_type, 16#0F#),
      3376 => to_slv(opcode_type, 16#0C#),
      3377 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#06#),
      3393 => to_slv(opcode_type, 16#04#),
      3394 => to_slv(opcode_type, 16#05#),
      3395 => to_slv(opcode_type, 16#09#),
      3396 => to_slv(opcode_type, 16#0B#),
      3397 => to_slv(opcode_type, 16#1E#),
      3398 => to_slv(opcode_type, 16#07#),
      3399 => to_slv(opcode_type, 16#07#),
      3400 => to_slv(opcode_type, 16#06#),
      3401 => to_slv(opcode_type, 16#5D#),
      3402 => to_slv(opcode_type, 16#0B#),
      3403 => to_slv(opcode_type, 16#08#),
      3404 => to_slv(opcode_type, 16#0B#),
      3405 => to_slv(opcode_type, 16#0E#),
      3406 => to_slv(opcode_type, 16#05#),
      3407 => to_slv(opcode_type, 16#05#),
      3408 => to_slv(opcode_type, 16#0A#),
      3409 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#07#),
      3425 => to_slv(opcode_type, 16#08#),
      3426 => to_slv(opcode_type, 16#05#),
      3427 => to_slv(opcode_type, 16#04#),
      3428 => to_slv(opcode_type, 16#0F#),
      3429 => to_slv(opcode_type, 16#07#),
      3430 => to_slv(opcode_type, 16#02#),
      3431 => to_slv(opcode_type, 16#0E#),
      3432 => to_slv(opcode_type, 16#07#),
      3433 => to_slv(opcode_type, 16#0B#),
      3434 => to_slv(opcode_type, 16#0F#),
      3435 => to_slv(opcode_type, 16#07#),
      3436 => to_slv(opcode_type, 16#06#),
      3437 => to_slv(opcode_type, 16#05#),
      3438 => to_slv(opcode_type, 16#10#),
      3439 => to_slv(opcode_type, 16#15#),
      3440 => to_slv(opcode_type, 16#0F#),
      3441 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#06#),
      3457 => to_slv(opcode_type, 16#04#),
      3458 => to_slv(opcode_type, 16#03#),
      3459 => to_slv(opcode_type, 16#04#),
      3460 => to_slv(opcode_type, 16#0F#),
      3461 => to_slv(opcode_type, 16#09#),
      3462 => to_slv(opcode_type, 16#06#),
      3463 => to_slv(opcode_type, 16#02#),
      3464 => to_slv(opcode_type, 16#B9#),
      3465 => to_slv(opcode_type, 16#06#),
      3466 => to_slv(opcode_type, 16#0B#),
      3467 => to_slv(opcode_type, 16#0D#),
      3468 => to_slv(opcode_type, 16#08#),
      3469 => to_slv(opcode_type, 16#05#),
      3470 => to_slv(opcode_type, 16#0B#),
      3471 => to_slv(opcode_type, 16#01#),
      3472 => to_slv(opcode_type, 16#0B#),
      3473 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#06#),
      3489 => to_slv(opcode_type, 16#05#),
      3490 => to_slv(opcode_type, 16#03#),
      3491 => to_slv(opcode_type, 16#05#),
      3492 => to_slv(opcode_type, 16#0A#),
      3493 => to_slv(opcode_type, 16#06#),
      3494 => to_slv(opcode_type, 16#01#),
      3495 => to_slv(opcode_type, 16#06#),
      3496 => to_slv(opcode_type, 16#0C#),
      3497 => to_slv(opcode_type, 16#10#),
      3498 => to_slv(opcode_type, 16#08#),
      3499 => to_slv(opcode_type, 16#06#),
      3500 => to_slv(opcode_type, 16#0D#),
      3501 => to_slv(opcode_type, 16#0A#),
      3502 => to_slv(opcode_type, 16#08#),
      3503 => to_slv(opcode_type, 16#0C#),
      3504 => to_slv(opcode_type, 16#0C#),
      3505 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#07#),
      3521 => to_slv(opcode_type, 16#01#),
      3522 => to_slv(opcode_type, 16#08#),
      3523 => to_slv(opcode_type, 16#05#),
      3524 => to_slv(opcode_type, 16#0D#),
      3525 => to_slv(opcode_type, 16#02#),
      3526 => to_slv(opcode_type, 16#10#),
      3527 => to_slv(opcode_type, 16#06#),
      3528 => to_slv(opcode_type, 16#08#),
      3529 => to_slv(opcode_type, 16#04#),
      3530 => to_slv(opcode_type, 16#0B#),
      3531 => to_slv(opcode_type, 16#04#),
      3532 => to_slv(opcode_type, 16#0C#),
      3533 => to_slv(opcode_type, 16#01#),
      3534 => to_slv(opcode_type, 16#07#),
      3535 => to_slv(opcode_type, 16#0F#),
      3536 => to_slv(opcode_type, 16#0D#),
      3537 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#08#),
      3553 => to_slv(opcode_type, 16#01#),
      3554 => to_slv(opcode_type, 16#04#),
      3555 => to_slv(opcode_type, 16#02#),
      3556 => to_slv(opcode_type, 16#0F#),
      3557 => to_slv(opcode_type, 16#09#),
      3558 => to_slv(opcode_type, 16#02#),
      3559 => to_slv(opcode_type, 16#09#),
      3560 => to_slv(opcode_type, 16#0E#),
      3561 => to_slv(opcode_type, 16#B4#),
      3562 => to_slv(opcode_type, 16#09#),
      3563 => to_slv(opcode_type, 16#06#),
      3564 => to_slv(opcode_type, 16#11#),
      3565 => to_slv(opcode_type, 16#0A#),
      3566 => to_slv(opcode_type, 16#06#),
      3567 => to_slv(opcode_type, 16#10#),
      3568 => to_slv(opcode_type, 16#0C#),
      3569 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#06#),
      3585 => to_slv(opcode_type, 16#07#),
      3586 => to_slv(opcode_type, 16#05#),
      3587 => to_slv(opcode_type, 16#02#),
      3588 => to_slv(opcode_type, 16#0E#),
      3589 => to_slv(opcode_type, 16#02#),
      3590 => to_slv(opcode_type, 16#02#),
      3591 => to_slv(opcode_type, 16#0B#),
      3592 => to_slv(opcode_type, 16#09#),
      3593 => to_slv(opcode_type, 16#01#),
      3594 => to_slv(opcode_type, 16#03#),
      3595 => to_slv(opcode_type, 16#5E#),
      3596 => to_slv(opcode_type, 16#09#),
      3597 => to_slv(opcode_type, 16#07#),
      3598 => to_slv(opcode_type, 16#0B#),
      3599 => to_slv(opcode_type, 16#0F#),
      3600 => to_slv(opcode_type, 16#0F#),
      3601 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#07#),
      3617 => to_slv(opcode_type, 16#05#),
      3618 => to_slv(opcode_type, 16#04#),
      3619 => to_slv(opcode_type, 16#01#),
      3620 => to_slv(opcode_type, 16#0F#),
      3621 => to_slv(opcode_type, 16#07#),
      3622 => to_slv(opcode_type, 16#09#),
      3623 => to_slv(opcode_type, 16#05#),
      3624 => to_slv(opcode_type, 16#10#),
      3625 => to_slv(opcode_type, 16#03#),
      3626 => to_slv(opcode_type, 16#E5#),
      3627 => to_slv(opcode_type, 16#07#),
      3628 => to_slv(opcode_type, 16#04#),
      3629 => to_slv(opcode_type, 16#10#),
      3630 => to_slv(opcode_type, 16#08#),
      3631 => to_slv(opcode_type, 16#0F#),
      3632 => to_slv(opcode_type, 16#11#),
      3633 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#08#),
      3649 => to_slv(opcode_type, 16#05#),
      3650 => to_slv(opcode_type, 16#06#),
      3651 => to_slv(opcode_type, 16#08#),
      3652 => to_slv(opcode_type, 16#0D#),
      3653 => to_slv(opcode_type, 16#0D#),
      3654 => to_slv(opcode_type, 16#09#),
      3655 => to_slv(opcode_type, 16#0A#),
      3656 => to_slv(opcode_type, 16#0A#),
      3657 => to_slv(opcode_type, 16#07#),
      3658 => to_slv(opcode_type, 16#05#),
      3659 => to_slv(opcode_type, 16#09#),
      3660 => to_slv(opcode_type, 16#0C#),
      3661 => to_slv(opcode_type, 16#11#),
      3662 => to_slv(opcode_type, 16#09#),
      3663 => to_slv(opcode_type, 16#11#),
      3664 => to_slv(opcode_type, 16#0C#),
      3665 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#09#),
      3681 => to_slv(opcode_type, 16#05#),
      3682 => to_slv(opcode_type, 16#01#),
      3683 => to_slv(opcode_type, 16#04#),
      3684 => to_slv(opcode_type, 16#0A#),
      3685 => to_slv(opcode_type, 16#08#),
      3686 => to_slv(opcode_type, 16#01#),
      3687 => to_slv(opcode_type, 16#07#),
      3688 => to_slv(opcode_type, 16#0C#),
      3689 => to_slv(opcode_type, 16#0F#),
      3690 => to_slv(opcode_type, 16#08#),
      3691 => to_slv(opcode_type, 16#07#),
      3692 => to_slv(opcode_type, 16#0D#),
      3693 => to_slv(opcode_type, 16#0A#),
      3694 => to_slv(opcode_type, 16#08#),
      3695 => to_slv(opcode_type, 16#0A#),
      3696 => to_slv(opcode_type, 16#9F#),
      3697 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#07#),
      3713 => to_slv(opcode_type, 16#04#),
      3714 => to_slv(opcode_type, 16#05#),
      3715 => to_slv(opcode_type, 16#05#),
      3716 => to_slv(opcode_type, 16#0C#),
      3717 => to_slv(opcode_type, 16#08#),
      3718 => to_slv(opcode_type, 16#05#),
      3719 => to_slv(opcode_type, 16#09#),
      3720 => to_slv(opcode_type, 16#0B#),
      3721 => to_slv(opcode_type, 16#0C#),
      3722 => to_slv(opcode_type, 16#06#),
      3723 => to_slv(opcode_type, 16#08#),
      3724 => to_slv(opcode_type, 16#0A#),
      3725 => to_slv(opcode_type, 16#0F#),
      3726 => to_slv(opcode_type, 16#09#),
      3727 => to_slv(opcode_type, 16#0C#),
      3728 => to_slv(opcode_type, 16#10#),
      3729 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#08#),
      3745 => to_slv(opcode_type, 16#04#),
      3746 => to_slv(opcode_type, 16#05#),
      3747 => to_slv(opcode_type, 16#08#),
      3748 => to_slv(opcode_type, 16#0F#),
      3749 => to_slv(opcode_type, 16#0B#),
      3750 => to_slv(opcode_type, 16#06#),
      3751 => to_slv(opcode_type, 16#09#),
      3752 => to_slv(opcode_type, 16#02#),
      3753 => to_slv(opcode_type, 16#0E#),
      3754 => to_slv(opcode_type, 16#02#),
      3755 => to_slv(opcode_type, 16#0D#),
      3756 => to_slv(opcode_type, 16#09#),
      3757 => to_slv(opcode_type, 16#09#),
      3758 => to_slv(opcode_type, 16#0E#),
      3759 => to_slv(opcode_type, 16#0A#),
      3760 => to_slv(opcode_type, 16#0B#),
      3761 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#06#),
      3777 => to_slv(opcode_type, 16#08#),
      3778 => to_slv(opcode_type, 16#01#),
      3779 => to_slv(opcode_type, 16#03#),
      3780 => to_slv(opcode_type, 16#10#),
      3781 => to_slv(opcode_type, 16#07#),
      3782 => to_slv(opcode_type, 16#05#),
      3783 => to_slv(opcode_type, 16#0E#),
      3784 => to_slv(opcode_type, 16#07#),
      3785 => to_slv(opcode_type, 16#0A#),
      3786 => to_slv(opcode_type, 16#0C#),
      3787 => to_slv(opcode_type, 16#03#),
      3788 => to_slv(opcode_type, 16#08#),
      3789 => to_slv(opcode_type, 16#07#),
      3790 => to_slv(opcode_type, 16#10#),
      3791 => to_slv(opcode_type, 16#0B#),
      3792 => to_slv(opcode_type, 16#0F#),
      3793 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#08#),
      3809 => to_slv(opcode_type, 16#09#),
      3810 => to_slv(opcode_type, 16#08#),
      3811 => to_slv(opcode_type, 16#09#),
      3812 => to_slv(opcode_type, 16#11#),
      3813 => to_slv(opcode_type, 16#0E#),
      3814 => to_slv(opcode_type, 16#01#),
      3815 => to_slv(opcode_type, 16#0F#),
      3816 => to_slv(opcode_type, 16#02#),
      3817 => to_slv(opcode_type, 16#01#),
      3818 => to_slv(opcode_type, 16#0F#),
      3819 => to_slv(opcode_type, 16#03#),
      3820 => to_slv(opcode_type, 16#06#),
      3821 => to_slv(opcode_type, 16#04#),
      3822 => to_slv(opcode_type, 16#0F#),
      3823 => to_slv(opcode_type, 16#05#),
      3824 => to_slv(opcode_type, 16#0D#),
      3825 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#09#),
      3841 => to_slv(opcode_type, 16#06#),
      3842 => to_slv(opcode_type, 16#08#),
      3843 => to_slv(opcode_type, 16#03#),
      3844 => to_slv(opcode_type, 16#0D#),
      3845 => to_slv(opcode_type, 16#06#),
      3846 => to_slv(opcode_type, 16#10#),
      3847 => to_slv(opcode_type, 16#0B#),
      3848 => to_slv(opcode_type, 16#07#),
      3849 => to_slv(opcode_type, 16#06#),
      3850 => to_slv(opcode_type, 16#0B#),
      3851 => to_slv(opcode_type, 16#0E#),
      3852 => to_slv(opcode_type, 16#08#),
      3853 => to_slv(opcode_type, 16#0F#),
      3854 => to_slv(opcode_type, 16#0C#),
      3855 => to_slv(opcode_type, 16#03#),
      3856 => to_slv(opcode_type, 16#0E#),
      3857 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#06#),
      3873 => to_slv(opcode_type, 16#09#),
      3874 => to_slv(opcode_type, 16#06#),
      3875 => to_slv(opcode_type, 16#09#),
      3876 => to_slv(opcode_type, 16#0E#),
      3877 => to_slv(opcode_type, 16#27#),
      3878 => to_slv(opcode_type, 16#02#),
      3879 => to_slv(opcode_type, 16#10#),
      3880 => to_slv(opcode_type, 16#02#),
      3881 => to_slv(opcode_type, 16#02#),
      3882 => to_slv(opcode_type, 16#0D#),
      3883 => to_slv(opcode_type, 16#04#),
      3884 => to_slv(opcode_type, 16#06#),
      3885 => to_slv(opcode_type, 16#05#),
      3886 => to_slv(opcode_type, 16#0F#),
      3887 => to_slv(opcode_type, 16#01#),
      3888 => to_slv(opcode_type, 16#0B#),
      3889 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#08#),
      3905 => to_slv(opcode_type, 16#01#),
      3906 => to_slv(opcode_type, 16#02#),
      3907 => to_slv(opcode_type, 16#08#),
      3908 => to_slv(opcode_type, 16#11#),
      3909 => to_slv(opcode_type, 16#0A#),
      3910 => to_slv(opcode_type, 16#08#),
      3911 => to_slv(opcode_type, 16#06#),
      3912 => to_slv(opcode_type, 16#03#),
      3913 => to_slv(opcode_type, 16#0A#),
      3914 => to_slv(opcode_type, 16#04#),
      3915 => to_slv(opcode_type, 16#11#),
      3916 => to_slv(opcode_type, 16#07#),
      3917 => to_slv(opcode_type, 16#05#),
      3918 => to_slv(opcode_type, 16#0F#),
      3919 => to_slv(opcode_type, 16#01#),
      3920 => to_slv(opcode_type, 16#0D#),
      3921 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#06#),
      3937 => to_slv(opcode_type, 16#09#),
      3938 => to_slv(opcode_type, 16#01#),
      3939 => to_slv(opcode_type, 16#06#),
      3940 => to_slv(opcode_type, 16#0B#),
      3941 => to_slv(opcode_type, 16#0E#),
      3942 => to_slv(opcode_type, 16#08#),
      3943 => to_slv(opcode_type, 16#04#),
      3944 => to_slv(opcode_type, 16#0B#),
      3945 => to_slv(opcode_type, 16#03#),
      3946 => to_slv(opcode_type, 16#0B#),
      3947 => to_slv(opcode_type, 16#09#),
      3948 => to_slv(opcode_type, 16#09#),
      3949 => to_slv(opcode_type, 16#01#),
      3950 => to_slv(opcode_type, 16#0C#),
      3951 => to_slv(opcode_type, 16#0B#),
      3952 => to_slv(opcode_type, 16#11#),
      3953 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#07#),
      3969 => to_slv(opcode_type, 16#04#),
      3970 => to_slv(opcode_type, 16#09#),
      3971 => to_slv(opcode_type, 16#09#),
      3972 => to_slv(opcode_type, 16#0F#),
      3973 => to_slv(opcode_type, 16#11#),
      3974 => to_slv(opcode_type, 16#03#),
      3975 => to_slv(opcode_type, 16#11#),
      3976 => to_slv(opcode_type, 16#06#),
      3977 => to_slv(opcode_type, 16#08#),
      3978 => to_slv(opcode_type, 16#09#),
      3979 => to_slv(opcode_type, 16#B6#),
      3980 => to_slv(opcode_type, 16#0D#),
      3981 => to_slv(opcode_type, 16#01#),
      3982 => to_slv(opcode_type, 16#0D#),
      3983 => to_slv(opcode_type, 16#05#),
      3984 => to_slv(opcode_type, 16#0F#),
      3985 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#07#),
      4001 => to_slv(opcode_type, 16#07#),
      4002 => to_slv(opcode_type, 16#06#),
      4003 => to_slv(opcode_type, 16#02#),
      4004 => to_slv(opcode_type, 16#10#),
      4005 => to_slv(opcode_type, 16#03#),
      4006 => to_slv(opcode_type, 16#0D#),
      4007 => to_slv(opcode_type, 16#03#),
      4008 => to_slv(opcode_type, 16#04#),
      4009 => to_slv(opcode_type, 16#0D#),
      4010 => to_slv(opcode_type, 16#03#),
      4011 => to_slv(opcode_type, 16#09#),
      4012 => to_slv(opcode_type, 16#06#),
      4013 => to_slv(opcode_type, 16#A3#),
      4014 => to_slv(opcode_type, 16#0E#),
      4015 => to_slv(opcode_type, 16#05#),
      4016 => to_slv(opcode_type, 16#0C#),
      4017 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#07#),
      4033 => to_slv(opcode_type, 16#01#),
      4034 => to_slv(opcode_type, 16#04#),
      4035 => to_slv(opcode_type, 16#03#),
      4036 => to_slv(opcode_type, 16#0F#),
      4037 => to_slv(opcode_type, 16#09#),
      4038 => to_slv(opcode_type, 16#01#),
      4039 => to_slv(opcode_type, 16#08#),
      4040 => to_slv(opcode_type, 16#0B#),
      4041 => to_slv(opcode_type, 16#10#),
      4042 => to_slv(opcode_type, 16#08#),
      4043 => to_slv(opcode_type, 16#08#),
      4044 => to_slv(opcode_type, 16#0E#),
      4045 => to_slv(opcode_type, 16#11#),
      4046 => to_slv(opcode_type, 16#08#),
      4047 => to_slv(opcode_type, 16#0C#),
      4048 => to_slv(opcode_type, 16#0A#),
      4049 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#08#),
      4065 => to_slv(opcode_type, 16#01#),
      4066 => to_slv(opcode_type, 16#04#),
      4067 => to_slv(opcode_type, 16#05#),
      4068 => to_slv(opcode_type, 16#0D#),
      4069 => to_slv(opcode_type, 16#09#),
      4070 => to_slv(opcode_type, 16#06#),
      4071 => to_slv(opcode_type, 16#09#),
      4072 => to_slv(opcode_type, 16#0F#),
      4073 => to_slv(opcode_type, 16#0E#),
      4074 => to_slv(opcode_type, 16#08#),
      4075 => to_slv(opcode_type, 16#0C#),
      4076 => to_slv(opcode_type, 16#11#),
      4077 => to_slv(opcode_type, 16#07#),
      4078 => to_slv(opcode_type, 16#03#),
      4079 => to_slv(opcode_type, 16#7B#),
      4080 => to_slv(opcode_type, 16#11#),
      4081 to 4095 => (others => '0')
  ),

    -- Bin `18`...
    17 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#09#),
      1 => to_slv(opcode_type, 16#07#),
      2 => to_slv(opcode_type, 16#01#),
      3 => to_slv(opcode_type, 16#08#),
      4 => to_slv(opcode_type, 16#0E#),
      5 => to_slv(opcode_type, 16#11#),
      6 => to_slv(opcode_type, 16#01#),
      7 => to_slv(opcode_type, 16#04#),
      8 => to_slv(opcode_type, 16#0D#),
      9 => to_slv(opcode_type, 16#08#),
      10 => to_slv(opcode_type, 16#08#),
      11 => to_slv(opcode_type, 16#03#),
      12 => to_slv(opcode_type, 16#0F#),
      13 => to_slv(opcode_type, 16#05#),
      14 => to_slv(opcode_type, 16#0A#),
      15 => to_slv(opcode_type, 16#09#),
      16 => to_slv(opcode_type, 16#0C#),
      17 => to_slv(opcode_type, 16#0D#),
      18 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#08#),
      33 => to_slv(opcode_type, 16#09#),
      34 => to_slv(opcode_type, 16#02#),
      35 => to_slv(opcode_type, 16#01#),
      36 => to_slv(opcode_type, 16#10#),
      37 => to_slv(opcode_type, 16#08#),
      38 => to_slv(opcode_type, 16#09#),
      39 => to_slv(opcode_type, 16#0E#),
      40 => to_slv(opcode_type, 16#0E#),
      41 => to_slv(opcode_type, 16#01#),
      42 => to_slv(opcode_type, 16#0D#),
      43 => to_slv(opcode_type, 16#02#),
      44 => to_slv(opcode_type, 16#07#),
      45 => to_slv(opcode_type, 16#05#),
      46 => to_slv(opcode_type, 16#10#),
      47 => to_slv(opcode_type, 16#07#),
      48 => to_slv(opcode_type, 16#0A#),
      49 => to_slv(opcode_type, 16#11#),
      50 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#06#),
      65 => to_slv(opcode_type, 16#01#),
      66 => to_slv(opcode_type, 16#01#),
      67 => to_slv(opcode_type, 16#08#),
      68 => to_slv(opcode_type, 16#0C#),
      69 => to_slv(opcode_type, 16#10#),
      70 => to_slv(opcode_type, 16#08#),
      71 => to_slv(opcode_type, 16#02#),
      72 => to_slv(opcode_type, 16#09#),
      73 => to_slv(opcode_type, 16#11#),
      74 => to_slv(opcode_type, 16#8D#),
      75 => to_slv(opcode_type, 16#08#),
      76 => to_slv(opcode_type, 16#09#),
      77 => to_slv(opcode_type, 16#0A#),
      78 => to_slv(opcode_type, 16#0D#),
      79 => to_slv(opcode_type, 16#07#),
      80 => to_slv(opcode_type, 16#11#),
      81 => to_slv(opcode_type, 16#0B#),
      82 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#06#),
      97 => to_slv(opcode_type, 16#08#),
      98 => to_slv(opcode_type, 16#01#),
      99 => to_slv(opcode_type, 16#03#),
      100 => to_slv(opcode_type, 16#0D#),
      101 => to_slv(opcode_type, 16#06#),
      102 => to_slv(opcode_type, 16#03#),
      103 => to_slv(opcode_type, 16#2E#),
      104 => to_slv(opcode_type, 16#05#),
      105 => to_slv(opcode_type, 16#0A#),
      106 => to_slv(opcode_type, 16#04#),
      107 => to_slv(opcode_type, 16#07#),
      108 => to_slv(opcode_type, 16#08#),
      109 => to_slv(opcode_type, 16#0A#),
      110 => to_slv(opcode_type, 16#0B#),
      111 => to_slv(opcode_type, 16#09#),
      112 => to_slv(opcode_type, 16#0F#),
      113 => to_slv(opcode_type, 16#0A#),
      114 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#06#),
      129 => to_slv(opcode_type, 16#05#),
      130 => to_slv(opcode_type, 16#06#),
      131 => to_slv(opcode_type, 16#04#),
      132 => to_slv(opcode_type, 16#0B#),
      133 => to_slv(opcode_type, 16#08#),
      134 => to_slv(opcode_type, 16#11#),
      135 => to_slv(opcode_type, 16#10#),
      136 => to_slv(opcode_type, 16#08#),
      137 => to_slv(opcode_type, 16#04#),
      138 => to_slv(opcode_type, 16#01#),
      139 => to_slv(opcode_type, 16#0A#),
      140 => to_slv(opcode_type, 16#06#),
      141 => to_slv(opcode_type, 16#04#),
      142 => to_slv(opcode_type, 16#10#),
      143 => to_slv(opcode_type, 16#06#),
      144 => to_slv(opcode_type, 16#0F#),
      145 => to_slv(opcode_type, 16#0C#),
      146 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#09#),
      161 => to_slv(opcode_type, 16#03#),
      162 => to_slv(opcode_type, 16#01#),
      163 => to_slv(opcode_type, 16#09#),
      164 => to_slv(opcode_type, 16#0E#),
      165 => to_slv(opcode_type, 16#0A#),
      166 => to_slv(opcode_type, 16#07#),
      167 => to_slv(opcode_type, 16#09#),
      168 => to_slv(opcode_type, 16#01#),
      169 => to_slv(opcode_type, 16#DC#),
      170 => to_slv(opcode_type, 16#08#),
      171 => to_slv(opcode_type, 16#0B#),
      172 => to_slv(opcode_type, 16#D2#),
      173 => to_slv(opcode_type, 16#09#),
      174 => to_slv(opcode_type, 16#03#),
      175 => to_slv(opcode_type, 16#0A#),
      176 => to_slv(opcode_type, 16#03#),
      177 => to_slv(opcode_type, 16#0A#),
      178 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#08#),
      193 => to_slv(opcode_type, 16#03#),
      194 => to_slv(opcode_type, 16#05#),
      195 => to_slv(opcode_type, 16#09#),
      196 => to_slv(opcode_type, 16#79#),
      197 => to_slv(opcode_type, 16#0B#),
      198 => to_slv(opcode_type, 16#08#),
      199 => to_slv(opcode_type, 16#01#),
      200 => to_slv(opcode_type, 16#07#),
      201 => to_slv(opcode_type, 16#0F#),
      202 => to_slv(opcode_type, 16#0C#),
      203 => to_slv(opcode_type, 16#09#),
      204 => to_slv(opcode_type, 16#08#),
      205 => to_slv(opcode_type, 16#10#),
      206 => to_slv(opcode_type, 16#66#),
      207 => to_slv(opcode_type, 16#08#),
      208 => to_slv(opcode_type, 16#0B#),
      209 => to_slv(opcode_type, 16#10#),
      210 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#07#),
      225 => to_slv(opcode_type, 16#07#),
      226 => to_slv(opcode_type, 16#09#),
      227 => to_slv(opcode_type, 16#01#),
      228 => to_slv(opcode_type, 16#0B#),
      229 => to_slv(opcode_type, 16#09#),
      230 => to_slv(opcode_type, 16#0E#),
      231 => to_slv(opcode_type, 16#11#),
      232 => to_slv(opcode_type, 16#03#),
      233 => to_slv(opcode_type, 16#06#),
      234 => to_slv(opcode_type, 16#0C#),
      235 => to_slv(opcode_type, 16#11#),
      236 => to_slv(opcode_type, 16#07#),
      237 => to_slv(opcode_type, 16#09#),
      238 => to_slv(opcode_type, 16#04#),
      239 => to_slv(opcode_type, 16#0E#),
      240 => to_slv(opcode_type, 16#1A#),
      241 => to_slv(opcode_type, 16#10#),
      242 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#07#),
      257 => to_slv(opcode_type, 16#07#),
      258 => to_slv(opcode_type, 16#04#),
      259 => to_slv(opcode_type, 16#01#),
      260 => to_slv(opcode_type, 16#0E#),
      261 => to_slv(opcode_type, 16#03#),
      262 => to_slv(opcode_type, 16#01#),
      263 => to_slv(opcode_type, 16#0E#),
      264 => to_slv(opcode_type, 16#06#),
      265 => to_slv(opcode_type, 16#06#),
      266 => to_slv(opcode_type, 16#07#),
      267 => to_slv(opcode_type, 16#10#),
      268 => to_slv(opcode_type, 16#11#),
      269 => to_slv(opcode_type, 16#06#),
      270 => to_slv(opcode_type, 16#11#),
      271 => to_slv(opcode_type, 16#0E#),
      272 => to_slv(opcode_type, 16#03#),
      273 => to_slv(opcode_type, 16#0E#),
      274 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#08#),
      290 => to_slv(opcode_type, 16#07#),
      291 => to_slv(opcode_type, 16#09#),
      292 => to_slv(opcode_type, 16#0E#),
      293 => to_slv(opcode_type, 16#94#),
      294 => to_slv(opcode_type, 16#05#),
      295 => to_slv(opcode_type, 16#11#),
      296 => to_slv(opcode_type, 16#09#),
      297 => to_slv(opcode_type, 16#08#),
      298 => to_slv(opcode_type, 16#11#),
      299 => to_slv(opcode_type, 16#0E#),
      300 => to_slv(opcode_type, 16#08#),
      301 => to_slv(opcode_type, 16#9D#),
      302 => to_slv(opcode_type, 16#B9#),
      303 => to_slv(opcode_type, 16#07#),
      304 => to_slv(opcode_type, 16#0B#),
      305 => to_slv(opcode_type, 16#0A#),
      306 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#09#),
      321 => to_slv(opcode_type, 16#04#),
      322 => to_slv(opcode_type, 16#07#),
      323 => to_slv(opcode_type, 16#02#),
      324 => to_slv(opcode_type, 16#0E#),
      325 => to_slv(opcode_type, 16#05#),
      326 => to_slv(opcode_type, 16#0A#),
      327 => to_slv(opcode_type, 16#07#),
      328 => to_slv(opcode_type, 16#04#),
      329 => to_slv(opcode_type, 16#08#),
      330 => to_slv(opcode_type, 16#10#),
      331 => to_slv(opcode_type, 16#0C#),
      332 => to_slv(opcode_type, 16#08#),
      333 => to_slv(opcode_type, 16#08#),
      334 => to_slv(opcode_type, 16#0B#),
      335 => to_slv(opcode_type, 16#FF#),
      336 => to_slv(opcode_type, 16#01#),
      337 => to_slv(opcode_type, 16#0A#),
      338 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#09#),
      353 => to_slv(opcode_type, 16#08#),
      354 => to_slv(opcode_type, 16#04#),
      355 => to_slv(opcode_type, 16#06#),
      356 => to_slv(opcode_type, 16#0E#),
      357 => to_slv(opcode_type, 16#4C#),
      358 => to_slv(opcode_type, 16#03#),
      359 => to_slv(opcode_type, 16#03#),
      360 => to_slv(opcode_type, 16#4A#),
      361 => to_slv(opcode_type, 16#08#),
      362 => to_slv(opcode_type, 16#08#),
      363 => to_slv(opcode_type, 16#07#),
      364 => to_slv(opcode_type, 16#10#),
      365 => to_slv(opcode_type, 16#0D#),
      366 => to_slv(opcode_type, 16#01#),
      367 => to_slv(opcode_type, 16#8D#),
      368 => to_slv(opcode_type, 16#04#),
      369 => to_slv(opcode_type, 16#0B#),
      370 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#09#),
      385 => to_slv(opcode_type, 16#08#),
      386 => to_slv(opcode_type, 16#01#),
      387 => to_slv(opcode_type, 16#01#),
      388 => to_slv(opcode_type, 16#0C#),
      389 => to_slv(opcode_type, 16#02#),
      390 => to_slv(opcode_type, 16#05#),
      391 => to_slv(opcode_type, 16#0E#),
      392 => to_slv(opcode_type, 16#08#),
      393 => to_slv(opcode_type, 16#03#),
      394 => to_slv(opcode_type, 16#02#),
      395 => to_slv(opcode_type, 16#0A#),
      396 => to_slv(opcode_type, 16#07#),
      397 => to_slv(opcode_type, 16#05#),
      398 => to_slv(opcode_type, 16#0B#),
      399 => to_slv(opcode_type, 16#06#),
      400 => to_slv(opcode_type, 16#10#),
      401 => to_slv(opcode_type, 16#0D#),
      402 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#06#),
      417 => to_slv(opcode_type, 16#09#),
      418 => to_slv(opcode_type, 16#03#),
      419 => to_slv(opcode_type, 16#04#),
      420 => to_slv(opcode_type, 16#10#),
      421 => to_slv(opcode_type, 16#06#),
      422 => to_slv(opcode_type, 16#05#),
      423 => to_slv(opcode_type, 16#0D#),
      424 => to_slv(opcode_type, 16#05#),
      425 => to_slv(opcode_type, 16#0C#),
      426 => to_slv(opcode_type, 16#08#),
      427 => to_slv(opcode_type, 16#02#),
      428 => to_slv(opcode_type, 16#02#),
      429 => to_slv(opcode_type, 16#0C#),
      430 => to_slv(opcode_type, 16#08#),
      431 => to_slv(opcode_type, 16#02#),
      432 => to_slv(opcode_type, 16#41#),
      433 => to_slv(opcode_type, 16#C1#),
      434 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#08#),
      449 => to_slv(opcode_type, 16#03#),
      450 => to_slv(opcode_type, 16#01#),
      451 => to_slv(opcode_type, 16#02#),
      452 => to_slv(opcode_type, 16#10#),
      453 => to_slv(opcode_type, 16#07#),
      454 => to_slv(opcode_type, 16#07#),
      455 => to_slv(opcode_type, 16#09#),
      456 => to_slv(opcode_type, 16#0E#),
      457 => to_slv(opcode_type, 16#0D#),
      458 => to_slv(opcode_type, 16#04#),
      459 => to_slv(opcode_type, 16#0B#),
      460 => to_slv(opcode_type, 16#09#),
      461 => to_slv(opcode_type, 16#09#),
      462 => to_slv(opcode_type, 16#0A#),
      463 => to_slv(opcode_type, 16#0F#),
      464 => to_slv(opcode_type, 16#04#),
      465 => to_slv(opcode_type, 16#10#),
      466 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#09#),
      481 => to_slv(opcode_type, 16#02#),
      482 => to_slv(opcode_type, 16#07#),
      483 => to_slv(opcode_type, 16#01#),
      484 => to_slv(opcode_type, 16#0A#),
      485 => to_slv(opcode_type, 16#03#),
      486 => to_slv(opcode_type, 16#0E#),
      487 => to_slv(opcode_type, 16#09#),
      488 => to_slv(opcode_type, 16#06#),
      489 => to_slv(opcode_type, 16#05#),
      490 => to_slv(opcode_type, 16#0B#),
      491 => to_slv(opcode_type, 16#08#),
      492 => to_slv(opcode_type, 16#F9#),
      493 => to_slv(opcode_type, 16#0E#),
      494 => to_slv(opcode_type, 16#02#),
      495 => to_slv(opcode_type, 16#06#),
      496 => to_slv(opcode_type, 16#11#),
      497 => to_slv(opcode_type, 16#11#),
      498 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#08#),
      513 => to_slv(opcode_type, 16#02#),
      514 => to_slv(opcode_type, 16#05#),
      515 => to_slv(opcode_type, 16#04#),
      516 => to_slv(opcode_type, 16#0E#),
      517 => to_slv(opcode_type, 16#07#),
      518 => to_slv(opcode_type, 16#09#),
      519 => to_slv(opcode_type, 16#06#),
      520 => to_slv(opcode_type, 16#0A#),
      521 => to_slv(opcode_type, 16#0C#),
      522 => to_slv(opcode_type, 16#08#),
      523 => to_slv(opcode_type, 16#7A#),
      524 => to_slv(opcode_type, 16#10#),
      525 => to_slv(opcode_type, 16#08#),
      526 => to_slv(opcode_type, 16#03#),
      527 => to_slv(opcode_type, 16#0E#),
      528 => to_slv(opcode_type, 16#01#),
      529 => to_slv(opcode_type, 16#1E#),
      530 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#09#),
      545 => to_slv(opcode_type, 16#02#),
      546 => to_slv(opcode_type, 16#04#),
      547 => to_slv(opcode_type, 16#02#),
      548 => to_slv(opcode_type, 16#90#),
      549 => to_slv(opcode_type, 16#06#),
      550 => to_slv(opcode_type, 16#06#),
      551 => to_slv(opcode_type, 16#07#),
      552 => to_slv(opcode_type, 16#0F#),
      553 => to_slv(opcode_type, 16#0B#),
      554 => to_slv(opcode_type, 16#07#),
      555 => to_slv(opcode_type, 16#0F#),
      556 => to_slv(opcode_type, 16#11#),
      557 => to_slv(opcode_type, 16#06#),
      558 => to_slv(opcode_type, 16#01#),
      559 => to_slv(opcode_type, 16#10#),
      560 => to_slv(opcode_type, 16#05#),
      561 => to_slv(opcode_type, 16#0F#),
      562 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#06#),
      577 => to_slv(opcode_type, 16#01#),
      578 => to_slv(opcode_type, 16#01#),
      579 => to_slv(opcode_type, 16#09#),
      580 => to_slv(opcode_type, 16#BD#),
      581 => to_slv(opcode_type, 16#10#),
      582 => to_slv(opcode_type, 16#07#),
      583 => to_slv(opcode_type, 16#01#),
      584 => to_slv(opcode_type, 16#06#),
      585 => to_slv(opcode_type, 16#0E#),
      586 => to_slv(opcode_type, 16#0C#),
      587 => to_slv(opcode_type, 16#09#),
      588 => to_slv(opcode_type, 16#08#),
      589 => to_slv(opcode_type, 16#10#),
      590 => to_slv(opcode_type, 16#E4#),
      591 => to_slv(opcode_type, 16#08#),
      592 => to_slv(opcode_type, 16#0F#),
      593 => to_slv(opcode_type, 16#0A#),
      594 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#08#),
      609 => to_slv(opcode_type, 16#06#),
      610 => to_slv(opcode_type, 16#02#),
      611 => to_slv(opcode_type, 16#05#),
      612 => to_slv(opcode_type, 16#0F#),
      613 => to_slv(opcode_type, 16#06#),
      614 => to_slv(opcode_type, 16#03#),
      615 => to_slv(opcode_type, 16#0A#),
      616 => to_slv(opcode_type, 16#07#),
      617 => to_slv(opcode_type, 16#56#),
      618 => to_slv(opcode_type, 16#F9#),
      619 => to_slv(opcode_type, 16#05#),
      620 => to_slv(opcode_type, 16#08#),
      621 => to_slv(opcode_type, 16#02#),
      622 => to_slv(opcode_type, 16#10#),
      623 => to_slv(opcode_type, 16#06#),
      624 => to_slv(opcode_type, 16#0F#),
      625 => to_slv(opcode_type, 16#CB#),
      626 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#08#),
      641 => to_slv(opcode_type, 16#05#),
      642 => to_slv(opcode_type, 16#06#),
      643 => to_slv(opcode_type, 16#09#),
      644 => to_slv(opcode_type, 16#0F#),
      645 => to_slv(opcode_type, 16#10#),
      646 => to_slv(opcode_type, 16#05#),
      647 => to_slv(opcode_type, 16#0F#),
      648 => to_slv(opcode_type, 16#07#),
      649 => to_slv(opcode_type, 16#08#),
      650 => to_slv(opcode_type, 16#03#),
      651 => to_slv(opcode_type, 16#0C#),
      652 => to_slv(opcode_type, 16#06#),
      653 => to_slv(opcode_type, 16#0E#),
      654 => to_slv(opcode_type, 16#0E#),
      655 => to_slv(opcode_type, 16#01#),
      656 => to_slv(opcode_type, 16#02#),
      657 => to_slv(opcode_type, 16#10#),
      658 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#09#),
      673 => to_slv(opcode_type, 16#01#),
      674 => to_slv(opcode_type, 16#09#),
      675 => to_slv(opcode_type, 16#03#),
      676 => to_slv(opcode_type, 16#0B#),
      677 => to_slv(opcode_type, 16#01#),
      678 => to_slv(opcode_type, 16#0A#),
      679 => to_slv(opcode_type, 16#06#),
      680 => to_slv(opcode_type, 16#07#),
      681 => to_slv(opcode_type, 16#03#),
      682 => to_slv(opcode_type, 16#0B#),
      683 => to_slv(opcode_type, 16#04#),
      684 => to_slv(opcode_type, 16#0C#),
      685 => to_slv(opcode_type, 16#07#),
      686 => to_slv(opcode_type, 16#02#),
      687 => to_slv(opcode_type, 16#0F#),
      688 => to_slv(opcode_type, 16#01#),
      689 => to_slv(opcode_type, 16#11#),
      690 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#07#),
      705 => to_slv(opcode_type, 16#06#),
      706 => to_slv(opcode_type, 16#08#),
      707 => to_slv(opcode_type, 16#09#),
      708 => to_slv(opcode_type, 16#11#),
      709 => to_slv(opcode_type, 16#9B#),
      710 => to_slv(opcode_type, 16#07#),
      711 => to_slv(opcode_type, 16#0C#),
      712 => to_slv(opcode_type, 16#0D#),
      713 => to_slv(opcode_type, 16#07#),
      714 => to_slv(opcode_type, 16#03#),
      715 => to_slv(opcode_type, 16#0E#),
      716 => to_slv(opcode_type, 16#08#),
      717 => to_slv(opcode_type, 16#0D#),
      718 => to_slv(opcode_type, 16#11#),
      719 => to_slv(opcode_type, 16#02#),
      720 => to_slv(opcode_type, 16#02#),
      721 => to_slv(opcode_type, 16#11#),
      722 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#09#),
      737 => to_slv(opcode_type, 16#09#),
      738 => to_slv(opcode_type, 16#02#),
      739 => to_slv(opcode_type, 16#07#),
      740 => to_slv(opcode_type, 16#0E#),
      741 => to_slv(opcode_type, 16#10#),
      742 => to_slv(opcode_type, 16#08#),
      743 => to_slv(opcode_type, 16#03#),
      744 => to_slv(opcode_type, 16#0C#),
      745 => to_slv(opcode_type, 16#01#),
      746 => to_slv(opcode_type, 16#0A#),
      747 => to_slv(opcode_type, 16#01#),
      748 => to_slv(opcode_type, 16#09#),
      749 => to_slv(opcode_type, 16#04#),
      750 => to_slv(opcode_type, 16#10#),
      751 => to_slv(opcode_type, 16#06#),
      752 => to_slv(opcode_type, 16#0D#),
      753 => to_slv(opcode_type, 16#0C#),
      754 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#09#),
      769 => to_slv(opcode_type, 16#06#),
      770 => to_slv(opcode_type, 16#05#),
      771 => to_slv(opcode_type, 16#03#),
      772 => to_slv(opcode_type, 16#0F#),
      773 => to_slv(opcode_type, 16#01#),
      774 => to_slv(opcode_type, 16#06#),
      775 => to_slv(opcode_type, 16#0F#),
      776 => to_slv(opcode_type, 16#11#),
      777 => to_slv(opcode_type, 16#06#),
      778 => to_slv(opcode_type, 16#02#),
      779 => to_slv(opcode_type, 16#05#),
      780 => to_slv(opcode_type, 16#0D#),
      781 => to_slv(opcode_type, 16#06#),
      782 => to_slv(opcode_type, 16#02#),
      783 => to_slv(opcode_type, 16#0D#),
      784 => to_slv(opcode_type, 16#04#),
      785 => to_slv(opcode_type, 16#10#),
      786 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#07#),
      801 => to_slv(opcode_type, 16#05#),
      802 => to_slv(opcode_type, 16#09#),
      803 => to_slv(opcode_type, 16#03#),
      804 => to_slv(opcode_type, 16#0A#),
      805 => to_slv(opcode_type, 16#07#),
      806 => to_slv(opcode_type, 16#6B#),
      807 => to_slv(opcode_type, 16#0B#),
      808 => to_slv(opcode_type, 16#08#),
      809 => to_slv(opcode_type, 16#05#),
      810 => to_slv(opcode_type, 16#08#),
      811 => to_slv(opcode_type, 16#0D#),
      812 => to_slv(opcode_type, 16#0A#),
      813 => to_slv(opcode_type, 16#06#),
      814 => to_slv(opcode_type, 16#01#),
      815 => to_slv(opcode_type, 16#0E#),
      816 => to_slv(opcode_type, 16#05#),
      817 => to_slv(opcode_type, 16#0A#),
      818 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#07#),
      833 => to_slv(opcode_type, 16#07#),
      834 => to_slv(opcode_type, 16#05#),
      835 => to_slv(opcode_type, 16#05#),
      836 => to_slv(opcode_type, 16#0B#),
      837 => to_slv(opcode_type, 16#01#),
      838 => to_slv(opcode_type, 16#09#),
      839 => to_slv(opcode_type, 16#0B#),
      840 => to_slv(opcode_type, 16#0D#),
      841 => to_slv(opcode_type, 16#09#),
      842 => to_slv(opcode_type, 16#04#),
      843 => to_slv(opcode_type, 16#06#),
      844 => to_slv(opcode_type, 16#B9#),
      845 => to_slv(opcode_type, 16#10#),
      846 => to_slv(opcode_type, 16#04#),
      847 => to_slv(opcode_type, 16#07#),
      848 => to_slv(opcode_type, 16#0D#),
      849 => to_slv(opcode_type, 16#11#),
      850 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#08#),
      865 => to_slv(opcode_type, 16#07#),
      866 => to_slv(opcode_type, 16#02#),
      867 => to_slv(opcode_type, 16#09#),
      868 => to_slv(opcode_type, 16#0F#),
      869 => to_slv(opcode_type, 16#0D#),
      870 => to_slv(opcode_type, 16#07#),
      871 => to_slv(opcode_type, 16#03#),
      872 => to_slv(opcode_type, 16#0C#),
      873 => to_slv(opcode_type, 16#08#),
      874 => to_slv(opcode_type, 16#0F#),
      875 => to_slv(opcode_type, 16#0C#),
      876 => to_slv(opcode_type, 16#05#),
      877 => to_slv(opcode_type, 16#08#),
      878 => to_slv(opcode_type, 16#03#),
      879 => to_slv(opcode_type, 16#61#),
      880 => to_slv(opcode_type, 16#05#),
      881 => to_slv(opcode_type, 16#0A#),
      882 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#04#),
      898 => to_slv(opcode_type, 16#06#),
      899 => to_slv(opcode_type, 16#05#),
      900 => to_slv(opcode_type, 16#0D#),
      901 => to_slv(opcode_type, 16#08#),
      902 => to_slv(opcode_type, 16#10#),
      903 => to_slv(opcode_type, 16#E9#),
      904 => to_slv(opcode_type, 16#07#),
      905 => to_slv(opcode_type, 16#05#),
      906 => to_slv(opcode_type, 16#06#),
      907 => to_slv(opcode_type, 16#0F#),
      908 => to_slv(opcode_type, 16#0E#),
      909 => to_slv(opcode_type, 16#08#),
      910 => to_slv(opcode_type, 16#05#),
      911 => to_slv(opcode_type, 16#0D#),
      912 => to_slv(opcode_type, 16#03#),
      913 => to_slv(opcode_type, 16#0A#),
      914 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#06#),
      929 => to_slv(opcode_type, 16#03#),
      930 => to_slv(opcode_type, 16#05#),
      931 => to_slv(opcode_type, 16#04#),
      932 => to_slv(opcode_type, 16#11#),
      933 => to_slv(opcode_type, 16#07#),
      934 => to_slv(opcode_type, 16#07#),
      935 => to_slv(opcode_type, 16#07#),
      936 => to_slv(opcode_type, 16#0A#),
      937 => to_slv(opcode_type, 16#79#),
      938 => to_slv(opcode_type, 16#05#),
      939 => to_slv(opcode_type, 16#19#),
      940 => to_slv(opcode_type, 16#08#),
      941 => to_slv(opcode_type, 16#05#),
      942 => to_slv(opcode_type, 16#0C#),
      943 => to_slv(opcode_type, 16#08#),
      944 => to_slv(opcode_type, 16#0C#),
      945 => to_slv(opcode_type, 16#0B#),
      946 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#06#),
      961 => to_slv(opcode_type, 16#03#),
      962 => to_slv(opcode_type, 16#02#),
      963 => to_slv(opcode_type, 16#05#),
      964 => to_slv(opcode_type, 16#1D#),
      965 => to_slv(opcode_type, 16#09#),
      966 => to_slv(opcode_type, 16#08#),
      967 => to_slv(opcode_type, 16#06#),
      968 => to_slv(opcode_type, 16#0F#),
      969 => to_slv(opcode_type, 16#0F#),
      970 => to_slv(opcode_type, 16#09#),
      971 => to_slv(opcode_type, 16#11#),
      972 => to_slv(opcode_type, 16#0A#),
      973 => to_slv(opcode_type, 16#06#),
      974 => to_slv(opcode_type, 16#02#),
      975 => to_slv(opcode_type, 16#0A#),
      976 => to_slv(opcode_type, 16#03#),
      977 => to_slv(opcode_type, 16#0F#),
      978 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#06#),
      993 => to_slv(opcode_type, 16#09#),
      994 => to_slv(opcode_type, 16#07#),
      995 => to_slv(opcode_type, 16#08#),
      996 => to_slv(opcode_type, 16#10#),
      997 => to_slv(opcode_type, 16#11#),
      998 => to_slv(opcode_type, 16#06#),
      999 => to_slv(opcode_type, 16#10#),
      1000 => to_slv(opcode_type, 16#0C#),
      1001 => to_slv(opcode_type, 16#03#),
      1002 => to_slv(opcode_type, 16#09#),
      1003 => to_slv(opcode_type, 16#0D#),
      1004 => to_slv(opcode_type, 16#AE#),
      1005 => to_slv(opcode_type, 16#07#),
      1006 => to_slv(opcode_type, 16#04#),
      1007 => to_slv(opcode_type, 16#01#),
      1008 => to_slv(opcode_type, 16#11#),
      1009 => to_slv(opcode_type, 16#0D#),
      1010 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#09#),
      1025 => to_slv(opcode_type, 16#09#),
      1026 => to_slv(opcode_type, 16#06#),
      1027 => to_slv(opcode_type, 16#03#),
      1028 => to_slv(opcode_type, 16#0F#),
      1029 => to_slv(opcode_type, 16#09#),
      1030 => to_slv(opcode_type, 16#0B#),
      1031 => to_slv(opcode_type, 16#11#),
      1032 => to_slv(opcode_type, 16#09#),
      1033 => to_slv(opcode_type, 16#07#),
      1034 => to_slv(opcode_type, 16#0A#),
      1035 => to_slv(opcode_type, 16#10#),
      1036 => to_slv(opcode_type, 16#03#),
      1037 => to_slv(opcode_type, 16#10#),
      1038 => to_slv(opcode_type, 16#09#),
      1039 => to_slv(opcode_type, 16#04#),
      1040 => to_slv(opcode_type, 16#F3#),
      1041 => to_slv(opcode_type, 16#0A#),
      1042 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#07#),
      1057 => to_slv(opcode_type, 16#09#),
      1058 => to_slv(opcode_type, 16#09#),
      1059 => to_slv(opcode_type, 16#08#),
      1060 => to_slv(opcode_type, 16#0D#),
      1061 => to_slv(opcode_type, 16#11#),
      1062 => to_slv(opcode_type, 16#05#),
      1063 => to_slv(opcode_type, 16#0A#),
      1064 => to_slv(opcode_type, 16#02#),
      1065 => to_slv(opcode_type, 16#06#),
      1066 => to_slv(opcode_type, 16#0A#),
      1067 => to_slv(opcode_type, 16#0C#),
      1068 => to_slv(opcode_type, 16#09#),
      1069 => to_slv(opcode_type, 16#06#),
      1070 => to_slv(opcode_type, 16#04#),
      1071 => to_slv(opcode_type, 16#0A#),
      1072 => to_slv(opcode_type, 16#0A#),
      1073 => to_slv(opcode_type, 16#0D#),
      1074 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#09#),
      1089 => to_slv(opcode_type, 16#03#),
      1090 => to_slv(opcode_type, 16#04#),
      1091 => to_slv(opcode_type, 16#01#),
      1092 => to_slv(opcode_type, 16#26#),
      1093 => to_slv(opcode_type, 16#06#),
      1094 => to_slv(opcode_type, 16#08#),
      1095 => to_slv(opcode_type, 16#06#),
      1096 => to_slv(opcode_type, 16#10#),
      1097 => to_slv(opcode_type, 16#0A#),
      1098 => to_slv(opcode_type, 16#09#),
      1099 => to_slv(opcode_type, 16#0F#),
      1100 => to_slv(opcode_type, 16#D7#),
      1101 => to_slv(opcode_type, 16#09#),
      1102 => to_slv(opcode_type, 16#09#),
      1103 => to_slv(opcode_type, 16#0C#),
      1104 => to_slv(opcode_type, 16#11#),
      1105 => to_slv(opcode_type, 16#10#),
      1106 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#06#),
      1121 => to_slv(opcode_type, 16#06#),
      1122 => to_slv(opcode_type, 16#06#),
      1123 => to_slv(opcode_type, 16#07#),
      1124 => to_slv(opcode_type, 16#0B#),
      1125 => to_slv(opcode_type, 16#0C#),
      1126 => to_slv(opcode_type, 16#07#),
      1127 => to_slv(opcode_type, 16#33#),
      1128 => to_slv(opcode_type, 16#10#),
      1129 => to_slv(opcode_type, 16#06#),
      1130 => to_slv(opcode_type, 16#03#),
      1131 => to_slv(opcode_type, 16#11#),
      1132 => to_slv(opcode_type, 16#08#),
      1133 => to_slv(opcode_type, 16#0E#),
      1134 => to_slv(opcode_type, 16#11#),
      1135 => to_slv(opcode_type, 16#02#),
      1136 => to_slv(opcode_type, 16#03#),
      1137 => to_slv(opcode_type, 16#0D#),
      1138 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#06#),
      1153 => to_slv(opcode_type, 16#02#),
      1154 => to_slv(opcode_type, 16#08#),
      1155 => to_slv(opcode_type, 16#06#),
      1156 => to_slv(opcode_type, 16#0C#),
      1157 => to_slv(opcode_type, 16#0A#),
      1158 => to_slv(opcode_type, 16#04#),
      1159 => to_slv(opcode_type, 16#11#),
      1160 => to_slv(opcode_type, 16#08#),
      1161 => to_slv(opcode_type, 16#04#),
      1162 => to_slv(opcode_type, 16#09#),
      1163 => to_slv(opcode_type, 16#0D#),
      1164 => to_slv(opcode_type, 16#0E#),
      1165 => to_slv(opcode_type, 16#06#),
      1166 => to_slv(opcode_type, 16#05#),
      1167 => to_slv(opcode_type, 16#0C#),
      1168 => to_slv(opcode_type, 16#05#),
      1169 => to_slv(opcode_type, 16#0C#),
      1170 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#07#),
      1185 => to_slv(opcode_type, 16#09#),
      1186 => to_slv(opcode_type, 16#04#),
      1187 => to_slv(opcode_type, 16#04#),
      1188 => to_slv(opcode_type, 16#0C#),
      1189 => to_slv(opcode_type, 16#09#),
      1190 => to_slv(opcode_type, 16#02#),
      1191 => to_slv(opcode_type, 16#D3#),
      1192 => to_slv(opcode_type, 16#03#),
      1193 => to_slv(opcode_type, 16#10#),
      1194 => to_slv(opcode_type, 16#07#),
      1195 => to_slv(opcode_type, 16#07#),
      1196 => to_slv(opcode_type, 16#01#),
      1197 => to_slv(opcode_type, 16#11#),
      1198 => to_slv(opcode_type, 16#02#),
      1199 => to_slv(opcode_type, 16#0A#),
      1200 => to_slv(opcode_type, 16#01#),
      1201 => to_slv(opcode_type, 16#0D#),
      1202 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#08#),
      1217 => to_slv(opcode_type, 16#01#),
      1218 => to_slv(opcode_type, 16#08#),
      1219 => to_slv(opcode_type, 16#03#),
      1220 => to_slv(opcode_type, 16#31#),
      1221 => to_slv(opcode_type, 16#03#),
      1222 => to_slv(opcode_type, 16#0E#),
      1223 => to_slv(opcode_type, 16#08#),
      1224 => to_slv(opcode_type, 16#06#),
      1225 => to_slv(opcode_type, 16#02#),
      1226 => to_slv(opcode_type, 16#0E#),
      1227 => to_slv(opcode_type, 16#01#),
      1228 => to_slv(opcode_type, 16#0F#),
      1229 => to_slv(opcode_type, 16#09#),
      1230 => to_slv(opcode_type, 16#04#),
      1231 => to_slv(opcode_type, 16#0C#),
      1232 => to_slv(opcode_type, 16#05#),
      1233 => to_slv(opcode_type, 16#0F#),
      1234 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#06#),
      1249 => to_slv(opcode_type, 16#01#),
      1250 => to_slv(opcode_type, 16#09#),
      1251 => to_slv(opcode_type, 16#08#),
      1252 => to_slv(opcode_type, 16#0A#),
      1253 => to_slv(opcode_type, 16#0D#),
      1254 => to_slv(opcode_type, 16#04#),
      1255 => to_slv(opcode_type, 16#0C#),
      1256 => to_slv(opcode_type, 16#08#),
      1257 => to_slv(opcode_type, 16#08#),
      1258 => to_slv(opcode_type, 16#02#),
      1259 => to_slv(opcode_type, 16#5C#),
      1260 => to_slv(opcode_type, 16#05#),
      1261 => to_slv(opcode_type, 16#0A#),
      1262 => to_slv(opcode_type, 16#01#),
      1263 => to_slv(opcode_type, 16#09#),
      1264 => to_slv(opcode_type, 16#0A#),
      1265 => to_slv(opcode_type, 16#0C#),
      1266 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#08#),
      1282 => to_slv(opcode_type, 16#06#),
      1283 => to_slv(opcode_type, 16#02#),
      1284 => to_slv(opcode_type, 16#0B#),
      1285 => to_slv(opcode_type, 16#02#),
      1286 => to_slv(opcode_type, 16#0F#),
      1287 => to_slv(opcode_type, 16#02#),
      1288 => to_slv(opcode_type, 16#01#),
      1289 => to_slv(opcode_type, 16#0A#),
      1290 => to_slv(opcode_type, 16#06#),
      1291 => to_slv(opcode_type, 16#06#),
      1292 => to_slv(opcode_type, 16#08#),
      1293 => to_slv(opcode_type, 16#0E#),
      1294 => to_slv(opcode_type, 16#0F#),
      1295 => to_slv(opcode_type, 16#05#),
      1296 => to_slv(opcode_type, 16#0F#),
      1297 => to_slv(opcode_type, 16#0C#),
      1298 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#07#),
      1313 => to_slv(opcode_type, 16#03#),
      1314 => to_slv(opcode_type, 16#06#),
      1315 => to_slv(opcode_type, 16#02#),
      1316 => to_slv(opcode_type, 16#0A#),
      1317 => to_slv(opcode_type, 16#01#),
      1318 => to_slv(opcode_type, 16#0F#),
      1319 => to_slv(opcode_type, 16#09#),
      1320 => to_slv(opcode_type, 16#09#),
      1321 => to_slv(opcode_type, 16#09#),
      1322 => to_slv(opcode_type, 16#0F#),
      1323 => to_slv(opcode_type, 16#0A#),
      1324 => to_slv(opcode_type, 16#04#),
      1325 => to_slv(opcode_type, 16#0F#),
      1326 => to_slv(opcode_type, 16#07#),
      1327 => to_slv(opcode_type, 16#03#),
      1328 => to_slv(opcode_type, 16#0C#),
      1329 => to_slv(opcode_type, 16#0D#),
      1330 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#09#),
      1345 => to_slv(opcode_type, 16#04#),
      1346 => to_slv(opcode_type, 16#07#),
      1347 => to_slv(opcode_type, 16#04#),
      1348 => to_slv(opcode_type, 16#10#),
      1349 => to_slv(opcode_type, 16#02#),
      1350 => to_slv(opcode_type, 16#0D#),
      1351 => to_slv(opcode_type, 16#07#),
      1352 => to_slv(opcode_type, 16#01#),
      1353 => to_slv(opcode_type, 16#02#),
      1354 => to_slv(opcode_type, 16#0E#),
      1355 => to_slv(opcode_type, 16#08#),
      1356 => to_slv(opcode_type, 16#09#),
      1357 => to_slv(opcode_type, 16#10#),
      1358 => to_slv(opcode_type, 16#10#),
      1359 => to_slv(opcode_type, 16#09#),
      1360 => to_slv(opcode_type, 16#11#),
      1361 => to_slv(opcode_type, 16#0B#),
      1362 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#09#),
      1377 => to_slv(opcode_type, 16#09#),
      1378 => to_slv(opcode_type, 16#02#),
      1379 => to_slv(opcode_type, 16#01#),
      1380 => to_slv(opcode_type, 16#0E#),
      1381 => to_slv(opcode_type, 16#07#),
      1382 => to_slv(opcode_type, 16#04#),
      1383 => to_slv(opcode_type, 16#0E#),
      1384 => to_slv(opcode_type, 16#04#),
      1385 => to_slv(opcode_type, 16#11#),
      1386 => to_slv(opcode_type, 16#03#),
      1387 => to_slv(opcode_type, 16#08#),
      1388 => to_slv(opcode_type, 16#09#),
      1389 => to_slv(opcode_type, 16#0A#),
      1390 => to_slv(opcode_type, 16#0D#),
      1391 => to_slv(opcode_type, 16#07#),
      1392 => to_slv(opcode_type, 16#F8#),
      1393 => to_slv(opcode_type, 16#11#),
      1394 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#07#),
      1409 => to_slv(opcode_type, 16#06#),
      1410 => to_slv(opcode_type, 16#01#),
      1411 => to_slv(opcode_type, 16#04#),
      1412 => to_slv(opcode_type, 16#0F#),
      1413 => to_slv(opcode_type, 16#03#),
      1414 => to_slv(opcode_type, 16#05#),
      1415 => to_slv(opcode_type, 16#0E#),
      1416 => to_slv(opcode_type, 16#07#),
      1417 => to_slv(opcode_type, 16#01#),
      1418 => to_slv(opcode_type, 16#09#),
      1419 => to_slv(opcode_type, 16#11#),
      1420 => to_slv(opcode_type, 16#0C#),
      1421 => to_slv(opcode_type, 16#09#),
      1422 => to_slv(opcode_type, 16#01#),
      1423 => to_slv(opcode_type, 16#11#),
      1424 => to_slv(opcode_type, 16#05#),
      1425 => to_slv(opcode_type, 16#0A#),
      1426 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#09#),
      1441 => to_slv(opcode_type, 16#04#),
      1442 => to_slv(opcode_type, 16#08#),
      1443 => to_slv(opcode_type, 16#06#),
      1444 => to_slv(opcode_type, 16#0E#),
      1445 => to_slv(opcode_type, 16#0B#),
      1446 => to_slv(opcode_type, 16#01#),
      1447 => to_slv(opcode_type, 16#0B#),
      1448 => to_slv(opcode_type, 16#08#),
      1449 => to_slv(opcode_type, 16#05#),
      1450 => to_slv(opcode_type, 16#02#),
      1451 => to_slv(opcode_type, 16#0E#),
      1452 => to_slv(opcode_type, 16#08#),
      1453 => to_slv(opcode_type, 16#04#),
      1454 => to_slv(opcode_type, 16#0E#),
      1455 => to_slv(opcode_type, 16#08#),
      1456 => to_slv(opcode_type, 16#0F#),
      1457 => to_slv(opcode_type, 16#0A#),
      1458 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#07#),
      1473 => to_slv(opcode_type, 16#01#),
      1474 => to_slv(opcode_type, 16#09#),
      1475 => to_slv(opcode_type, 16#03#),
      1476 => to_slv(opcode_type, 16#0A#),
      1477 => to_slv(opcode_type, 16#02#),
      1478 => to_slv(opcode_type, 16#10#),
      1479 => to_slv(opcode_type, 16#07#),
      1480 => to_slv(opcode_type, 16#05#),
      1481 => to_slv(opcode_type, 16#01#),
      1482 => to_slv(opcode_type, 16#10#),
      1483 => to_slv(opcode_type, 16#08#),
      1484 => to_slv(opcode_type, 16#06#),
      1485 => to_slv(opcode_type, 16#0D#),
      1486 => to_slv(opcode_type, 16#10#),
      1487 => to_slv(opcode_type, 16#06#),
      1488 => to_slv(opcode_type, 16#0A#),
      1489 => to_slv(opcode_type, 16#11#),
      1490 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#08#),
      1505 => to_slv(opcode_type, 16#07#),
      1506 => to_slv(opcode_type, 16#03#),
      1507 => to_slv(opcode_type, 16#09#),
      1508 => to_slv(opcode_type, 16#26#),
      1509 => to_slv(opcode_type, 16#0B#),
      1510 => to_slv(opcode_type, 16#02#),
      1511 => to_slv(opcode_type, 16#08#),
      1512 => to_slv(opcode_type, 16#73#),
      1513 => to_slv(opcode_type, 16#0C#),
      1514 => to_slv(opcode_type, 16#09#),
      1515 => to_slv(opcode_type, 16#06#),
      1516 => to_slv(opcode_type, 16#08#),
      1517 => to_slv(opcode_type, 16#0F#),
      1518 => to_slv(opcode_type, 16#0C#),
      1519 => to_slv(opcode_type, 16#02#),
      1520 => to_slv(opcode_type, 16#0C#),
      1521 => to_slv(opcode_type, 16#11#),
      1522 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#07#),
      1537 => to_slv(opcode_type, 16#04#),
      1538 => to_slv(opcode_type, 16#09#),
      1539 => to_slv(opcode_type, 16#06#),
      1540 => to_slv(opcode_type, 16#11#),
      1541 => to_slv(opcode_type, 16#0B#),
      1542 => to_slv(opcode_type, 16#07#),
      1543 => to_slv(opcode_type, 16#0C#),
      1544 => to_slv(opcode_type, 16#0E#),
      1545 => to_slv(opcode_type, 16#07#),
      1546 => to_slv(opcode_type, 16#05#),
      1547 => to_slv(opcode_type, 16#05#),
      1548 => to_slv(opcode_type, 16#11#),
      1549 => to_slv(opcode_type, 16#09#),
      1550 => to_slv(opcode_type, 16#04#),
      1551 => to_slv(opcode_type, 16#0B#),
      1552 => to_slv(opcode_type, 16#01#),
      1553 => to_slv(opcode_type, 16#0A#),
      1554 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#09#),
      1569 => to_slv(opcode_type, 16#02#),
      1570 => to_slv(opcode_type, 16#05#),
      1571 => to_slv(opcode_type, 16#07#),
      1572 => to_slv(opcode_type, 16#10#),
      1573 => to_slv(opcode_type, 16#0F#),
      1574 => to_slv(opcode_type, 16#08#),
      1575 => to_slv(opcode_type, 16#01#),
      1576 => to_slv(opcode_type, 16#09#),
      1577 => to_slv(opcode_type, 16#11#),
      1578 => to_slv(opcode_type, 16#0E#),
      1579 => to_slv(opcode_type, 16#09#),
      1580 => to_slv(opcode_type, 16#07#),
      1581 => to_slv(opcode_type, 16#10#),
      1582 => to_slv(opcode_type, 16#10#),
      1583 => to_slv(opcode_type, 16#07#),
      1584 => to_slv(opcode_type, 16#0C#),
      1585 => to_slv(opcode_type, 16#0E#),
      1586 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#02#),
      1602 => to_slv(opcode_type, 16#06#),
      1603 => to_slv(opcode_type, 16#07#),
      1604 => to_slv(opcode_type, 16#0C#),
      1605 => to_slv(opcode_type, 16#0B#),
      1606 => to_slv(opcode_type, 16#08#),
      1607 => to_slv(opcode_type, 16#0B#),
      1608 => to_slv(opcode_type, 16#0F#),
      1609 => to_slv(opcode_type, 16#09#),
      1610 => to_slv(opcode_type, 16#06#),
      1611 => to_slv(opcode_type, 16#01#),
      1612 => to_slv(opcode_type, 16#0F#),
      1613 => to_slv(opcode_type, 16#09#),
      1614 => to_slv(opcode_type, 16#0A#),
      1615 => to_slv(opcode_type, 16#0A#),
      1616 => to_slv(opcode_type, 16#02#),
      1617 => to_slv(opcode_type, 16#11#),
      1618 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#09#),
      1633 => to_slv(opcode_type, 16#09#),
      1634 => to_slv(opcode_type, 16#07#),
      1635 => to_slv(opcode_type, 16#05#),
      1636 => to_slv(opcode_type, 16#11#),
      1637 => to_slv(opcode_type, 16#04#),
      1638 => to_slv(opcode_type, 16#11#),
      1639 => to_slv(opcode_type, 16#04#),
      1640 => to_slv(opcode_type, 16#04#),
      1641 => to_slv(opcode_type, 16#0D#),
      1642 => to_slv(opcode_type, 16#05#),
      1643 => to_slv(opcode_type, 16#08#),
      1644 => to_slv(opcode_type, 16#07#),
      1645 => to_slv(opcode_type, 16#0D#),
      1646 => to_slv(opcode_type, 16#0A#),
      1647 => to_slv(opcode_type, 16#08#),
      1648 => to_slv(opcode_type, 16#3A#),
      1649 => to_slv(opcode_type, 16#0A#),
      1650 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#07#),
      1665 => to_slv(opcode_type, 16#05#),
      1666 => to_slv(opcode_type, 16#06#),
      1667 => to_slv(opcode_type, 16#02#),
      1668 => to_slv(opcode_type, 16#0D#),
      1669 => to_slv(opcode_type, 16#07#),
      1670 => to_slv(opcode_type, 16#11#),
      1671 => to_slv(opcode_type, 16#D7#),
      1672 => to_slv(opcode_type, 16#07#),
      1673 => to_slv(opcode_type, 16#05#),
      1674 => to_slv(opcode_type, 16#07#),
      1675 => to_slv(opcode_type, 16#10#),
      1676 => to_slv(opcode_type, 16#11#),
      1677 => to_slv(opcode_type, 16#07#),
      1678 => to_slv(opcode_type, 16#09#),
      1679 => to_slv(opcode_type, 16#11#),
      1680 => to_slv(opcode_type, 16#10#),
      1681 => to_slv(opcode_type, 16#7F#),
      1682 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#08#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#05#),
      1699 => to_slv(opcode_type, 16#01#),
      1700 => to_slv(opcode_type, 16#0D#),
      1701 => to_slv(opcode_type, 16#09#),
      1702 => to_slv(opcode_type, 16#08#),
      1703 => to_slv(opcode_type, 16#F2#),
      1704 => to_slv(opcode_type, 16#0A#),
      1705 => to_slv(opcode_type, 16#09#),
      1706 => to_slv(opcode_type, 16#0F#),
      1707 => to_slv(opcode_type, 16#11#),
      1708 => to_slv(opcode_type, 16#06#),
      1709 => to_slv(opcode_type, 16#02#),
      1710 => to_slv(opcode_type, 16#08#),
      1711 => to_slv(opcode_type, 16#0E#),
      1712 => to_slv(opcode_type, 16#11#),
      1713 => to_slv(opcode_type, 16#0E#),
      1714 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#08#),
      1729 => to_slv(opcode_type, 16#04#),
      1730 => to_slv(opcode_type, 16#05#),
      1731 => to_slv(opcode_type, 16#01#),
      1732 => to_slv(opcode_type, 16#10#),
      1733 => to_slv(opcode_type, 16#07#),
      1734 => to_slv(opcode_type, 16#06#),
      1735 => to_slv(opcode_type, 16#06#),
      1736 => to_slv(opcode_type, 16#0F#),
      1737 => to_slv(opcode_type, 16#0E#),
      1738 => to_slv(opcode_type, 16#01#),
      1739 => to_slv(opcode_type, 16#0F#),
      1740 => to_slv(opcode_type, 16#07#),
      1741 => to_slv(opcode_type, 16#04#),
      1742 => to_slv(opcode_type, 16#0D#),
      1743 => to_slv(opcode_type, 16#09#),
      1744 => to_slv(opcode_type, 16#0D#),
      1745 => to_slv(opcode_type, 16#CB#),
      1746 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#06#),
      1761 => to_slv(opcode_type, 16#09#),
      1762 => to_slv(opcode_type, 16#03#),
      1763 => to_slv(opcode_type, 16#02#),
      1764 => to_slv(opcode_type, 16#81#),
      1765 => to_slv(opcode_type, 16#05#),
      1766 => to_slv(opcode_type, 16#08#),
      1767 => to_slv(opcode_type, 16#10#),
      1768 => to_slv(opcode_type, 16#0B#),
      1769 => to_slv(opcode_type, 16#08#),
      1770 => to_slv(opcode_type, 16#05#),
      1771 => to_slv(opcode_type, 16#05#),
      1772 => to_slv(opcode_type, 16#10#),
      1773 => to_slv(opcode_type, 16#09#),
      1774 => to_slv(opcode_type, 16#03#),
      1775 => to_slv(opcode_type, 16#10#),
      1776 => to_slv(opcode_type, 16#05#),
      1777 => to_slv(opcode_type, 16#0F#),
      1778 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#08#),
      1793 => to_slv(opcode_type, 16#04#),
      1794 => to_slv(opcode_type, 16#08#),
      1795 => to_slv(opcode_type, 16#02#),
      1796 => to_slv(opcode_type, 16#0C#),
      1797 => to_slv(opcode_type, 16#09#),
      1798 => to_slv(opcode_type, 16#11#),
      1799 => to_slv(opcode_type, 16#0B#),
      1800 => to_slv(opcode_type, 16#06#),
      1801 => to_slv(opcode_type, 16#07#),
      1802 => to_slv(opcode_type, 16#07#),
      1803 => to_slv(opcode_type, 16#1B#),
      1804 => to_slv(opcode_type, 16#0C#),
      1805 => to_slv(opcode_type, 16#04#),
      1806 => to_slv(opcode_type, 16#0F#),
      1807 => to_slv(opcode_type, 16#07#),
      1808 => to_slv(opcode_type, 16#0C#),
      1809 => to_slv(opcode_type, 16#0E#),
      1810 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#06#),
      1825 => to_slv(opcode_type, 16#01#),
      1826 => to_slv(opcode_type, 16#05#),
      1827 => to_slv(opcode_type, 16#02#),
      1828 => to_slv(opcode_type, 16#0C#),
      1829 => to_slv(opcode_type, 16#09#),
      1830 => to_slv(opcode_type, 16#08#),
      1831 => to_slv(opcode_type, 16#05#),
      1832 => to_slv(opcode_type, 16#0B#),
      1833 => to_slv(opcode_type, 16#04#),
      1834 => to_slv(opcode_type, 16#0F#),
      1835 => to_slv(opcode_type, 16#09#),
      1836 => to_slv(opcode_type, 16#09#),
      1837 => to_slv(opcode_type, 16#0F#),
      1838 => to_slv(opcode_type, 16#0A#),
      1839 => to_slv(opcode_type, 16#06#),
      1840 => to_slv(opcode_type, 16#0C#),
      1841 => to_slv(opcode_type, 16#0D#),
      1842 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#08#),
      1857 => to_slv(opcode_type, 16#09#),
      1858 => to_slv(opcode_type, 16#08#),
      1859 => to_slv(opcode_type, 16#07#),
      1860 => to_slv(opcode_type, 16#10#),
      1861 => to_slv(opcode_type, 16#10#),
      1862 => to_slv(opcode_type, 16#04#),
      1863 => to_slv(opcode_type, 16#10#),
      1864 => to_slv(opcode_type, 16#05#),
      1865 => to_slv(opcode_type, 16#03#),
      1866 => to_slv(opcode_type, 16#0B#),
      1867 => to_slv(opcode_type, 16#01#),
      1868 => to_slv(opcode_type, 16#08#),
      1869 => to_slv(opcode_type, 16#04#),
      1870 => to_slv(opcode_type, 16#11#),
      1871 => to_slv(opcode_type, 16#06#),
      1872 => to_slv(opcode_type, 16#37#),
      1873 => to_slv(opcode_type, 16#0C#),
      1874 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#06#),
      1890 => to_slv(opcode_type, 16#09#),
      1891 => to_slv(opcode_type, 16#08#),
      1892 => to_slv(opcode_type, 16#0A#),
      1893 => to_slv(opcode_type, 16#0B#),
      1894 => to_slv(opcode_type, 16#07#),
      1895 => to_slv(opcode_type, 16#0C#),
      1896 => to_slv(opcode_type, 16#0F#),
      1897 => to_slv(opcode_type, 16#08#),
      1898 => to_slv(opcode_type, 16#02#),
      1899 => to_slv(opcode_type, 16#10#),
      1900 => to_slv(opcode_type, 16#08#),
      1901 => to_slv(opcode_type, 16#0B#),
      1902 => to_slv(opcode_type, 16#0C#),
      1903 => to_slv(opcode_type, 16#09#),
      1904 => to_slv(opcode_type, 16#83#),
      1905 => to_slv(opcode_type, 16#0A#),
      1906 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#08#),
      1921 => to_slv(opcode_type, 16#03#),
      1922 => to_slv(opcode_type, 16#03#),
      1923 => to_slv(opcode_type, 16#07#),
      1924 => to_slv(opcode_type, 16#0A#),
      1925 => to_slv(opcode_type, 16#10#),
      1926 => to_slv(opcode_type, 16#06#),
      1927 => to_slv(opcode_type, 16#08#),
      1928 => to_slv(opcode_type, 16#09#),
      1929 => to_slv(opcode_type, 16#0C#),
      1930 => to_slv(opcode_type, 16#0C#),
      1931 => to_slv(opcode_type, 16#08#),
      1932 => to_slv(opcode_type, 16#0C#),
      1933 => to_slv(opcode_type, 16#0B#),
      1934 => to_slv(opcode_type, 16#03#),
      1935 => to_slv(opcode_type, 16#07#),
      1936 => to_slv(opcode_type, 16#0C#),
      1937 => to_slv(opcode_type, 16#0D#),
      1938 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#07#),
      1953 => to_slv(opcode_type, 16#05#),
      1954 => to_slv(opcode_type, 16#01#),
      1955 => to_slv(opcode_type, 16#02#),
      1956 => to_slv(opcode_type, 16#62#),
      1957 => to_slv(opcode_type, 16#09#),
      1958 => to_slv(opcode_type, 16#08#),
      1959 => to_slv(opcode_type, 16#06#),
      1960 => to_slv(opcode_type, 16#0F#),
      1961 => to_slv(opcode_type, 16#0E#),
      1962 => to_slv(opcode_type, 16#09#),
      1963 => to_slv(opcode_type, 16#10#),
      1964 => to_slv(opcode_type, 16#11#),
      1965 => to_slv(opcode_type, 16#06#),
      1966 => to_slv(opcode_type, 16#01#),
      1967 => to_slv(opcode_type, 16#0B#),
      1968 => to_slv(opcode_type, 16#02#),
      1969 => to_slv(opcode_type, 16#0C#),
      1970 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#08#),
      1985 => to_slv(opcode_type, 16#07#),
      1986 => to_slv(opcode_type, 16#03#),
      1987 => to_slv(opcode_type, 16#09#),
      1988 => to_slv(opcode_type, 16#0F#),
      1989 => to_slv(opcode_type, 16#0A#),
      1990 => to_slv(opcode_type, 16#09#),
      1991 => to_slv(opcode_type, 16#07#),
      1992 => to_slv(opcode_type, 16#0F#),
      1993 => to_slv(opcode_type, 16#0E#),
      1994 => to_slv(opcode_type, 16#05#),
      1995 => to_slv(opcode_type, 16#0A#),
      1996 => to_slv(opcode_type, 16#04#),
      1997 => to_slv(opcode_type, 16#07#),
      1998 => to_slv(opcode_type, 16#03#),
      1999 => to_slv(opcode_type, 16#0C#),
      2000 => to_slv(opcode_type, 16#01#),
      2001 => to_slv(opcode_type, 16#0E#),
      2002 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#08#),
      2017 => to_slv(opcode_type, 16#09#),
      2018 => to_slv(opcode_type, 16#01#),
      2019 => to_slv(opcode_type, 16#01#),
      2020 => to_slv(opcode_type, 16#0F#),
      2021 => to_slv(opcode_type, 16#09#),
      2022 => to_slv(opcode_type, 16#04#),
      2023 => to_slv(opcode_type, 16#3F#),
      2024 => to_slv(opcode_type, 16#04#),
      2025 => to_slv(opcode_type, 16#0F#),
      2026 => to_slv(opcode_type, 16#06#),
      2027 => to_slv(opcode_type, 16#02#),
      2028 => to_slv(opcode_type, 16#05#),
      2029 => to_slv(opcode_type, 16#0D#),
      2030 => to_slv(opcode_type, 16#09#),
      2031 => to_slv(opcode_type, 16#03#),
      2032 => to_slv(opcode_type, 16#0E#),
      2033 => to_slv(opcode_type, 16#0E#),
      2034 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#07#),
      2049 => to_slv(opcode_type, 16#04#),
      2050 => to_slv(opcode_type, 16#05#),
      2051 => to_slv(opcode_type, 16#05#),
      2052 => to_slv(opcode_type, 16#0D#),
      2053 => to_slv(opcode_type, 16#08#),
      2054 => to_slv(opcode_type, 16#09#),
      2055 => to_slv(opcode_type, 16#08#),
      2056 => to_slv(opcode_type, 16#0F#),
      2057 => to_slv(opcode_type, 16#11#),
      2058 => to_slv(opcode_type, 16#09#),
      2059 => to_slv(opcode_type, 16#0A#),
      2060 => to_slv(opcode_type, 16#0A#),
      2061 => to_slv(opcode_type, 16#08#),
      2062 => to_slv(opcode_type, 16#06#),
      2063 => to_slv(opcode_type, 16#0D#),
      2064 => to_slv(opcode_type, 16#10#),
      2065 => to_slv(opcode_type, 16#0F#),
      2066 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#07#),
      2081 => to_slv(opcode_type, 16#04#),
      2082 => to_slv(opcode_type, 16#08#),
      2083 => to_slv(opcode_type, 16#03#),
      2084 => to_slv(opcode_type, 16#0E#),
      2085 => to_slv(opcode_type, 16#04#),
      2086 => to_slv(opcode_type, 16#3B#),
      2087 => to_slv(opcode_type, 16#07#),
      2088 => to_slv(opcode_type, 16#03#),
      2089 => to_slv(opcode_type, 16#02#),
      2090 => to_slv(opcode_type, 16#0E#),
      2091 => to_slv(opcode_type, 16#09#),
      2092 => to_slv(opcode_type, 16#07#),
      2093 => to_slv(opcode_type, 16#11#),
      2094 => to_slv(opcode_type, 16#0E#),
      2095 => to_slv(opcode_type, 16#07#),
      2096 => to_slv(opcode_type, 16#2B#),
      2097 => to_slv(opcode_type, 16#0A#),
      2098 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#08#),
      2113 => to_slv(opcode_type, 16#05#),
      2114 => to_slv(opcode_type, 16#09#),
      2115 => to_slv(opcode_type, 16#07#),
      2116 => to_slv(opcode_type, 16#0E#),
      2117 => to_slv(opcode_type, 16#0B#),
      2118 => to_slv(opcode_type, 16#01#),
      2119 => to_slv(opcode_type, 16#10#),
      2120 => to_slv(opcode_type, 16#06#),
      2121 => to_slv(opcode_type, 16#08#),
      2122 => to_slv(opcode_type, 16#04#),
      2123 => to_slv(opcode_type, 16#74#),
      2124 => to_slv(opcode_type, 16#06#),
      2125 => to_slv(opcode_type, 16#10#),
      2126 => to_slv(opcode_type, 16#0A#),
      2127 => to_slv(opcode_type, 16#09#),
      2128 => to_slv(opcode_type, 16#0B#),
      2129 => to_slv(opcode_type, 16#0B#),
      2130 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#02#),
      2146 => to_slv(opcode_type, 16#05#),
      2147 => to_slv(opcode_type, 16#01#),
      2148 => to_slv(opcode_type, 16#1B#),
      2149 => to_slv(opcode_type, 16#08#),
      2150 => to_slv(opcode_type, 16#09#),
      2151 => to_slv(opcode_type, 16#08#),
      2152 => to_slv(opcode_type, 16#0B#),
      2153 => to_slv(opcode_type, 16#0E#),
      2154 => to_slv(opcode_type, 16#05#),
      2155 => to_slv(opcode_type, 16#0E#),
      2156 => to_slv(opcode_type, 16#07#),
      2157 => to_slv(opcode_type, 16#02#),
      2158 => to_slv(opcode_type, 16#0B#),
      2159 => to_slv(opcode_type, 16#09#),
      2160 => to_slv(opcode_type, 16#0E#),
      2161 => to_slv(opcode_type, 16#0D#),
      2162 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#08#),
      2177 => to_slv(opcode_type, 16#05#),
      2178 => to_slv(opcode_type, 16#09#),
      2179 => to_slv(opcode_type, 16#04#),
      2180 => to_slv(opcode_type, 16#FD#),
      2181 => to_slv(opcode_type, 16#07#),
      2182 => to_slv(opcode_type, 16#0D#),
      2183 => to_slv(opcode_type, 16#11#),
      2184 => to_slv(opcode_type, 16#08#),
      2185 => to_slv(opcode_type, 16#01#),
      2186 => to_slv(opcode_type, 16#09#),
      2187 => to_slv(opcode_type, 16#0B#),
      2188 => to_slv(opcode_type, 16#10#),
      2189 => to_slv(opcode_type, 16#07#),
      2190 => to_slv(opcode_type, 16#09#),
      2191 => to_slv(opcode_type, 16#0B#),
      2192 => to_slv(opcode_type, 16#4A#),
      2193 => to_slv(opcode_type, 16#0E#),
      2194 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#07#),
      2209 => to_slv(opcode_type, 16#01#),
      2210 => to_slv(opcode_type, 16#06#),
      2211 => to_slv(opcode_type, 16#05#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#07#),
      2214 => to_slv(opcode_type, 16#11#),
      2215 => to_slv(opcode_type, 16#0B#),
      2216 => to_slv(opcode_type, 16#07#),
      2217 => to_slv(opcode_type, 16#03#),
      2218 => to_slv(opcode_type, 16#02#),
      2219 => to_slv(opcode_type, 16#0F#),
      2220 => to_slv(opcode_type, 16#08#),
      2221 => to_slv(opcode_type, 16#01#),
      2222 => to_slv(opcode_type, 16#0F#),
      2223 => to_slv(opcode_type, 16#06#),
      2224 => to_slv(opcode_type, 16#0C#),
      2225 => to_slv(opcode_type, 16#11#),
      2226 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#05#),
      2242 => to_slv(opcode_type, 16#09#),
      2243 => to_slv(opcode_type, 16#02#),
      2244 => to_slv(opcode_type, 16#10#),
      2245 => to_slv(opcode_type, 16#01#),
      2246 => to_slv(opcode_type, 16#0E#),
      2247 => to_slv(opcode_type, 16#07#),
      2248 => to_slv(opcode_type, 16#01#),
      2249 => to_slv(opcode_type, 16#07#),
      2250 => to_slv(opcode_type, 16#0D#),
      2251 => to_slv(opcode_type, 16#0A#),
      2252 => to_slv(opcode_type, 16#06#),
      2253 => to_slv(opcode_type, 16#03#),
      2254 => to_slv(opcode_type, 16#10#),
      2255 => to_slv(opcode_type, 16#06#),
      2256 => to_slv(opcode_type, 16#0F#),
      2257 => to_slv(opcode_type, 16#0D#),
      2258 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#09#),
      2273 => to_slv(opcode_type, 16#01#),
      2274 => to_slv(opcode_type, 16#01#),
      2275 => to_slv(opcode_type, 16#01#),
      2276 => to_slv(opcode_type, 16#10#),
      2277 => to_slv(opcode_type, 16#09#),
      2278 => to_slv(opcode_type, 16#06#),
      2279 => to_slv(opcode_type, 16#07#),
      2280 => to_slv(opcode_type, 16#0A#),
      2281 => to_slv(opcode_type, 16#0F#),
      2282 => to_slv(opcode_type, 16#08#),
      2283 => to_slv(opcode_type, 16#11#),
      2284 => to_slv(opcode_type, 16#0A#),
      2285 => to_slv(opcode_type, 16#06#),
      2286 => to_slv(opcode_type, 16#08#),
      2287 => to_slv(opcode_type, 16#A8#),
      2288 => to_slv(opcode_type, 16#0C#),
      2289 => to_slv(opcode_type, 16#0B#),
      2290 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#08#),
      2305 => to_slv(opcode_type, 16#08#),
      2306 => to_slv(opcode_type, 16#08#),
      2307 => to_slv(opcode_type, 16#07#),
      2308 => to_slv(opcode_type, 16#0C#),
      2309 => to_slv(opcode_type, 16#A2#),
      2310 => to_slv(opcode_type, 16#01#),
      2311 => to_slv(opcode_type, 16#10#),
      2312 => to_slv(opcode_type, 16#06#),
      2313 => to_slv(opcode_type, 16#01#),
      2314 => to_slv(opcode_type, 16#11#),
      2315 => to_slv(opcode_type, 16#02#),
      2316 => to_slv(opcode_type, 16#2E#),
      2317 => to_slv(opcode_type, 16#01#),
      2318 => to_slv(opcode_type, 16#06#),
      2319 => to_slv(opcode_type, 16#05#),
      2320 => to_slv(opcode_type, 16#F0#),
      2321 => to_slv(opcode_type, 16#0E#),
      2322 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#09#),
      2337 => to_slv(opcode_type, 16#05#),
      2338 => to_slv(opcode_type, 16#08#),
      2339 => to_slv(opcode_type, 16#06#),
      2340 => to_slv(opcode_type, 16#10#),
      2341 => to_slv(opcode_type, 16#0F#),
      2342 => to_slv(opcode_type, 16#08#),
      2343 => to_slv(opcode_type, 16#10#),
      2344 => to_slv(opcode_type, 16#10#),
      2345 => to_slv(opcode_type, 16#06#),
      2346 => to_slv(opcode_type, 16#07#),
      2347 => to_slv(opcode_type, 16#06#),
      2348 => to_slv(opcode_type, 16#11#),
      2349 => to_slv(opcode_type, 16#0B#),
      2350 => to_slv(opcode_type, 16#06#),
      2351 => to_slv(opcode_type, 16#11#),
      2352 => to_slv(opcode_type, 16#0C#),
      2353 => to_slv(opcode_type, 16#10#),
      2354 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#06#),
      2369 => to_slv(opcode_type, 16#01#),
      2370 => to_slv(opcode_type, 16#06#),
      2371 => to_slv(opcode_type, 16#09#),
      2372 => to_slv(opcode_type, 16#0C#),
      2373 => to_slv(opcode_type, 16#0C#),
      2374 => to_slv(opcode_type, 16#01#),
      2375 => to_slv(opcode_type, 16#DD#),
      2376 => to_slv(opcode_type, 16#06#),
      2377 => to_slv(opcode_type, 16#05#),
      2378 => to_slv(opcode_type, 16#05#),
      2379 => to_slv(opcode_type, 16#10#),
      2380 => to_slv(opcode_type, 16#08#),
      2381 => to_slv(opcode_type, 16#06#),
      2382 => to_slv(opcode_type, 16#2B#),
      2383 => to_slv(opcode_type, 16#0D#),
      2384 => to_slv(opcode_type, 16#03#),
      2385 => to_slv(opcode_type, 16#11#),
      2386 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#08#),
      2401 => to_slv(opcode_type, 16#03#),
      2402 => to_slv(opcode_type, 16#02#),
      2403 => to_slv(opcode_type, 16#01#),
      2404 => to_slv(opcode_type, 16#0D#),
      2405 => to_slv(opcode_type, 16#07#),
      2406 => to_slv(opcode_type, 16#08#),
      2407 => to_slv(opcode_type, 16#05#),
      2408 => to_slv(opcode_type, 16#0B#),
      2409 => to_slv(opcode_type, 16#06#),
      2410 => to_slv(opcode_type, 16#0D#),
      2411 => to_slv(opcode_type, 16#0D#),
      2412 => to_slv(opcode_type, 16#09#),
      2413 => to_slv(opcode_type, 16#09#),
      2414 => to_slv(opcode_type, 16#0A#),
      2415 => to_slv(opcode_type, 16#B4#),
      2416 => to_slv(opcode_type, 16#05#),
      2417 => to_slv(opcode_type, 16#0E#),
      2418 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#07#),
      2433 => to_slv(opcode_type, 16#07#),
      2434 => to_slv(opcode_type, 16#01#),
      2435 => to_slv(opcode_type, 16#08#),
      2436 => to_slv(opcode_type, 16#0B#),
      2437 => to_slv(opcode_type, 16#0B#),
      2438 => to_slv(opcode_type, 16#07#),
      2439 => to_slv(opcode_type, 16#02#),
      2440 => to_slv(opcode_type, 16#0E#),
      2441 => to_slv(opcode_type, 16#06#),
      2442 => to_slv(opcode_type, 16#11#),
      2443 => to_slv(opcode_type, 16#0A#),
      2444 => to_slv(opcode_type, 16#06#),
      2445 => to_slv(opcode_type, 16#05#),
      2446 => to_slv(opcode_type, 16#09#),
      2447 => to_slv(opcode_type, 16#B9#),
      2448 => to_slv(opcode_type, 16#0E#),
      2449 => to_slv(opcode_type, 16#11#),
      2450 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#09#),
      2465 => to_slv(opcode_type, 16#04#),
      2466 => to_slv(opcode_type, 16#02#),
      2467 => to_slv(opcode_type, 16#07#),
      2468 => to_slv(opcode_type, 16#10#),
      2469 => to_slv(opcode_type, 16#0C#),
      2470 => to_slv(opcode_type, 16#09#),
      2471 => to_slv(opcode_type, 16#03#),
      2472 => to_slv(opcode_type, 16#09#),
      2473 => to_slv(opcode_type, 16#0C#),
      2474 => to_slv(opcode_type, 16#0F#),
      2475 => to_slv(opcode_type, 16#06#),
      2476 => to_slv(opcode_type, 16#07#),
      2477 => to_slv(opcode_type, 16#0D#),
      2478 => to_slv(opcode_type, 16#0B#),
      2479 => to_slv(opcode_type, 16#09#),
      2480 => to_slv(opcode_type, 16#0C#),
      2481 => to_slv(opcode_type, 16#10#),
      2482 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#07#),
      2497 => to_slv(opcode_type, 16#02#),
      2498 => to_slv(opcode_type, 16#07#),
      2499 => to_slv(opcode_type, 16#07#),
      2500 => to_slv(opcode_type, 16#10#),
      2501 => to_slv(opcode_type, 16#10#),
      2502 => to_slv(opcode_type, 16#02#),
      2503 => to_slv(opcode_type, 16#0B#),
      2504 => to_slv(opcode_type, 16#09#),
      2505 => to_slv(opcode_type, 16#09#),
      2506 => to_slv(opcode_type, 16#03#),
      2507 => to_slv(opcode_type, 16#0D#),
      2508 => to_slv(opcode_type, 16#01#),
      2509 => to_slv(opcode_type, 16#8D#),
      2510 => to_slv(opcode_type, 16#02#),
      2511 => to_slv(opcode_type, 16#09#),
      2512 => to_slv(opcode_type, 16#0D#),
      2513 => to_slv(opcode_type, 16#0F#),
      2514 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#09#),
      2529 => to_slv(opcode_type, 16#09#),
      2530 => to_slv(opcode_type, 16#07#),
      2531 => to_slv(opcode_type, 16#02#),
      2532 => to_slv(opcode_type, 16#0D#),
      2533 => to_slv(opcode_type, 16#06#),
      2534 => to_slv(opcode_type, 16#11#),
      2535 => to_slv(opcode_type, 16#73#),
      2536 => to_slv(opcode_type, 16#01#),
      2537 => to_slv(opcode_type, 16#08#),
      2538 => to_slv(opcode_type, 16#0A#),
      2539 => to_slv(opcode_type, 16#0D#),
      2540 => to_slv(opcode_type, 16#02#),
      2541 => to_slv(opcode_type, 16#07#),
      2542 => to_slv(opcode_type, 16#06#),
      2543 => to_slv(opcode_type, 16#10#),
      2544 => to_slv(opcode_type, 16#0F#),
      2545 => to_slv(opcode_type, 16#0F#),
      2546 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#08#),
      2561 => to_slv(opcode_type, 16#03#),
      2562 => to_slv(opcode_type, 16#06#),
      2563 => to_slv(opcode_type, 16#03#),
      2564 => to_slv(opcode_type, 16#0E#),
      2565 => to_slv(opcode_type, 16#01#),
      2566 => to_slv(opcode_type, 16#0A#),
      2567 => to_slv(opcode_type, 16#08#),
      2568 => to_slv(opcode_type, 16#06#),
      2569 => to_slv(opcode_type, 16#07#),
      2570 => to_slv(opcode_type, 16#11#),
      2571 => to_slv(opcode_type, 16#10#),
      2572 => to_slv(opcode_type, 16#03#),
      2573 => to_slv(opcode_type, 16#58#),
      2574 => to_slv(opcode_type, 16#09#),
      2575 => to_slv(opcode_type, 16#01#),
      2576 => to_slv(opcode_type, 16#0B#),
      2577 => to_slv(opcode_type, 16#0F#),
      2578 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#07#),
      2593 => to_slv(opcode_type, 16#05#),
      2594 => to_slv(opcode_type, 16#09#),
      2595 => to_slv(opcode_type, 16#09#),
      2596 => to_slv(opcode_type, 16#0B#),
      2597 => to_slv(opcode_type, 16#0B#),
      2598 => to_slv(opcode_type, 16#07#),
      2599 => to_slv(opcode_type, 16#11#),
      2600 => to_slv(opcode_type, 16#0F#),
      2601 => to_slv(opcode_type, 16#08#),
      2602 => to_slv(opcode_type, 16#05#),
      2603 => to_slv(opcode_type, 16#08#),
      2604 => to_slv(opcode_type, 16#0C#),
      2605 => to_slv(opcode_type, 16#73#),
      2606 => to_slv(opcode_type, 16#08#),
      2607 => to_slv(opcode_type, 16#02#),
      2608 => to_slv(opcode_type, 16#0C#),
      2609 => to_slv(opcode_type, 16#0E#),
      2610 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#06#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#08#),
      2627 => to_slv(opcode_type, 16#06#),
      2628 => to_slv(opcode_type, 16#11#),
      2629 => to_slv(opcode_type, 16#0B#),
      2630 => to_slv(opcode_type, 16#06#),
      2631 => to_slv(opcode_type, 16#11#),
      2632 => to_slv(opcode_type, 16#0D#),
      2633 => to_slv(opcode_type, 16#05#),
      2634 => to_slv(opcode_type, 16#05#),
      2635 => to_slv(opcode_type, 16#10#),
      2636 => to_slv(opcode_type, 16#07#),
      2637 => to_slv(opcode_type, 16#03#),
      2638 => to_slv(opcode_type, 16#01#),
      2639 => to_slv(opcode_type, 16#11#),
      2640 => to_slv(opcode_type, 16#01#),
      2641 => to_slv(opcode_type, 16#11#),
      2642 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#06#),
      2657 => to_slv(opcode_type, 16#07#),
      2658 => to_slv(opcode_type, 16#07#),
      2659 => to_slv(opcode_type, 16#08#),
      2660 => to_slv(opcode_type, 16#0E#),
      2661 => to_slv(opcode_type, 16#0C#),
      2662 => to_slv(opcode_type, 16#06#),
      2663 => to_slv(opcode_type, 16#0F#),
      2664 => to_slv(opcode_type, 16#10#),
      2665 => to_slv(opcode_type, 16#09#),
      2666 => to_slv(opcode_type, 16#02#),
      2667 => to_slv(opcode_type, 16#0B#),
      2668 => to_slv(opcode_type, 16#08#),
      2669 => to_slv(opcode_type, 16#11#),
      2670 => to_slv(opcode_type, 16#6C#),
      2671 => to_slv(opcode_type, 16#01#),
      2672 => to_slv(opcode_type, 16#04#),
      2673 => to_slv(opcode_type, 16#0F#),
      2674 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#08#),
      2689 => to_slv(opcode_type, 16#03#),
      2690 => to_slv(opcode_type, 16#08#),
      2691 => to_slv(opcode_type, 16#02#),
      2692 => to_slv(opcode_type, 16#52#),
      2693 => to_slv(opcode_type, 16#04#),
      2694 => to_slv(opcode_type, 16#0F#),
      2695 => to_slv(opcode_type, 16#06#),
      2696 => to_slv(opcode_type, 16#01#),
      2697 => to_slv(opcode_type, 16#05#),
      2698 => to_slv(opcode_type, 16#11#),
      2699 => to_slv(opcode_type, 16#09#),
      2700 => to_slv(opcode_type, 16#09#),
      2701 => to_slv(opcode_type, 16#0F#),
      2702 => to_slv(opcode_type, 16#0F#),
      2703 => to_slv(opcode_type, 16#07#),
      2704 => to_slv(opcode_type, 16#10#),
      2705 => to_slv(opcode_type, 16#0F#),
      2706 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#06#),
      2721 => to_slv(opcode_type, 16#06#),
      2722 => to_slv(opcode_type, 16#07#),
      2723 => to_slv(opcode_type, 16#01#),
      2724 => to_slv(opcode_type, 16#11#),
      2725 => to_slv(opcode_type, 16#06#),
      2726 => to_slv(opcode_type, 16#0F#),
      2727 => to_slv(opcode_type, 16#0F#),
      2728 => to_slv(opcode_type, 16#06#),
      2729 => to_slv(opcode_type, 16#04#),
      2730 => to_slv(opcode_type, 16#0A#),
      2731 => to_slv(opcode_type, 16#01#),
      2732 => to_slv(opcode_type, 16#0A#),
      2733 => to_slv(opcode_type, 16#06#),
      2734 => to_slv(opcode_type, 16#02#),
      2735 => to_slv(opcode_type, 16#01#),
      2736 => to_slv(opcode_type, 16#11#),
      2737 => to_slv(opcode_type, 16#5D#),
      2738 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#07#),
      2753 => to_slv(opcode_type, 16#09#),
      2754 => to_slv(opcode_type, 16#03#),
      2755 => to_slv(opcode_type, 16#02#),
      2756 => to_slv(opcode_type, 16#0D#),
      2757 => to_slv(opcode_type, 16#09#),
      2758 => to_slv(opcode_type, 16#05#),
      2759 => to_slv(opcode_type, 16#0D#),
      2760 => to_slv(opcode_type, 16#02#),
      2761 => to_slv(opcode_type, 16#0E#),
      2762 => to_slv(opcode_type, 16#06#),
      2763 => to_slv(opcode_type, 16#05#),
      2764 => to_slv(opcode_type, 16#08#),
      2765 => to_slv(opcode_type, 16#0A#),
      2766 => to_slv(opcode_type, 16#0A#),
      2767 => to_slv(opcode_type, 16#08#),
      2768 => to_slv(opcode_type, 16#0F#),
      2769 => to_slv(opcode_type, 16#A0#),
      2770 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#07#),
      2785 => to_slv(opcode_type, 16#08#),
      2786 => to_slv(opcode_type, 16#03#),
      2787 => to_slv(opcode_type, 16#09#),
      2788 => to_slv(opcode_type, 16#0D#),
      2789 => to_slv(opcode_type, 16#0D#),
      2790 => to_slv(opcode_type, 16#08#),
      2791 => to_slv(opcode_type, 16#07#),
      2792 => to_slv(opcode_type, 16#0A#),
      2793 => to_slv(opcode_type, 16#0A#),
      2794 => to_slv(opcode_type, 16#06#),
      2795 => to_slv(opcode_type, 16#0A#),
      2796 => to_slv(opcode_type, 16#11#),
      2797 => to_slv(opcode_type, 16#03#),
      2798 => to_slv(opcode_type, 16#06#),
      2799 => to_slv(opcode_type, 16#03#),
      2800 => to_slv(opcode_type, 16#11#),
      2801 => to_slv(opcode_type, 16#0E#),
      2802 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#09#),
      2817 => to_slv(opcode_type, 16#01#),
      2818 => to_slv(opcode_type, 16#08#),
      2819 => to_slv(opcode_type, 16#03#),
      2820 => to_slv(opcode_type, 16#0B#),
      2821 => to_slv(opcode_type, 16#03#),
      2822 => to_slv(opcode_type, 16#11#),
      2823 => to_slv(opcode_type, 16#09#),
      2824 => to_slv(opcode_type, 16#09#),
      2825 => to_slv(opcode_type, 16#06#),
      2826 => to_slv(opcode_type, 16#0A#),
      2827 => to_slv(opcode_type, 16#0B#),
      2828 => to_slv(opcode_type, 16#06#),
      2829 => to_slv(opcode_type, 16#0E#),
      2830 => to_slv(opcode_type, 16#0E#),
      2831 => to_slv(opcode_type, 16#05#),
      2832 => to_slv(opcode_type, 16#02#),
      2833 => to_slv(opcode_type, 16#C2#),
      2834 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#06#),
      2849 => to_slv(opcode_type, 16#07#),
      2850 => to_slv(opcode_type, 16#08#),
      2851 => to_slv(opcode_type, 16#05#),
      2852 => to_slv(opcode_type, 16#10#),
      2853 => to_slv(opcode_type, 16#05#),
      2854 => to_slv(opcode_type, 16#0E#),
      2855 => to_slv(opcode_type, 16#05#),
      2856 => to_slv(opcode_type, 16#03#),
      2857 => to_slv(opcode_type, 16#0F#),
      2858 => to_slv(opcode_type, 16#09#),
      2859 => to_slv(opcode_type, 16#09#),
      2860 => to_slv(opcode_type, 16#09#),
      2861 => to_slv(opcode_type, 16#0C#),
      2862 => to_slv(opcode_type, 16#0E#),
      2863 => to_slv(opcode_type, 16#01#),
      2864 => to_slv(opcode_type, 16#0A#),
      2865 => to_slv(opcode_type, 16#0A#),
      2866 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#07#),
      2881 => to_slv(opcode_type, 16#05#),
      2882 => to_slv(opcode_type, 16#01#),
      2883 => to_slv(opcode_type, 16#02#),
      2884 => to_slv(opcode_type, 16#6D#),
      2885 => to_slv(opcode_type, 16#07#),
      2886 => to_slv(opcode_type, 16#09#),
      2887 => to_slv(opcode_type, 16#02#),
      2888 => to_slv(opcode_type, 16#0F#),
      2889 => to_slv(opcode_type, 16#05#),
      2890 => to_slv(opcode_type, 16#11#),
      2891 => to_slv(opcode_type, 16#08#),
      2892 => to_slv(opcode_type, 16#08#),
      2893 => to_slv(opcode_type, 16#10#),
      2894 => to_slv(opcode_type, 16#0B#),
      2895 => to_slv(opcode_type, 16#06#),
      2896 => to_slv(opcode_type, 16#0D#),
      2897 => to_slv(opcode_type, 16#0A#),
      2898 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#06#),
      2913 => to_slv(opcode_type, 16#04#),
      2914 => to_slv(opcode_type, 16#04#),
      2915 => to_slv(opcode_type, 16#01#),
      2916 => to_slv(opcode_type, 16#11#),
      2917 => to_slv(opcode_type, 16#08#),
      2918 => to_slv(opcode_type, 16#06#),
      2919 => to_slv(opcode_type, 16#03#),
      2920 => to_slv(opcode_type, 16#0F#),
      2921 => to_slv(opcode_type, 16#06#),
      2922 => to_slv(opcode_type, 16#0D#),
      2923 => to_slv(opcode_type, 16#10#),
      2924 => to_slv(opcode_type, 16#08#),
      2925 => to_slv(opcode_type, 16#02#),
      2926 => to_slv(opcode_type, 16#0F#),
      2927 => to_slv(opcode_type, 16#07#),
      2928 => to_slv(opcode_type, 16#0F#),
      2929 => to_slv(opcode_type, 16#0F#),
      2930 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#09#),
      2945 => to_slv(opcode_type, 16#06#),
      2946 => to_slv(opcode_type, 16#09#),
      2947 => to_slv(opcode_type, 16#02#),
      2948 => to_slv(opcode_type, 16#0A#),
      2949 => to_slv(opcode_type, 16#08#),
      2950 => to_slv(opcode_type, 16#11#),
      2951 => to_slv(opcode_type, 16#F1#),
      2952 => to_slv(opcode_type, 16#07#),
      2953 => to_slv(opcode_type, 16#05#),
      2954 => to_slv(opcode_type, 16#10#),
      2955 => to_slv(opcode_type, 16#04#),
      2956 => to_slv(opcode_type, 16#10#),
      2957 => to_slv(opcode_type, 16#03#),
      2958 => to_slv(opcode_type, 16#03#),
      2959 => to_slv(opcode_type, 16#07#),
      2960 => to_slv(opcode_type, 16#0F#),
      2961 => to_slv(opcode_type, 16#11#),
      2962 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#09#),
      2977 => to_slv(opcode_type, 16#04#),
      2978 => to_slv(opcode_type, 16#08#),
      2979 => to_slv(opcode_type, 16#01#),
      2980 => to_slv(opcode_type, 16#CB#),
      2981 => to_slv(opcode_type, 16#06#),
      2982 => to_slv(opcode_type, 16#92#),
      2983 => to_slv(opcode_type, 16#0F#),
      2984 => to_slv(opcode_type, 16#07#),
      2985 => to_slv(opcode_type, 16#07#),
      2986 => to_slv(opcode_type, 16#09#),
      2987 => to_slv(opcode_type, 16#0E#),
      2988 => to_slv(opcode_type, 16#0E#),
      2989 => to_slv(opcode_type, 16#04#),
      2990 => to_slv(opcode_type, 16#0A#),
      2991 => to_slv(opcode_type, 16#01#),
      2992 => to_slv(opcode_type, 16#04#),
      2993 => to_slv(opcode_type, 16#0D#),
      2994 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#08#),
      3009 => to_slv(opcode_type, 16#05#),
      3010 => to_slv(opcode_type, 16#05#),
      3011 => to_slv(opcode_type, 16#03#),
      3012 => to_slv(opcode_type, 16#0C#),
      3013 => to_slv(opcode_type, 16#07#),
      3014 => to_slv(opcode_type, 16#06#),
      3015 => to_slv(opcode_type, 16#08#),
      3016 => to_slv(opcode_type, 16#9E#),
      3017 => to_slv(opcode_type, 16#0E#),
      3018 => to_slv(opcode_type, 16#01#),
      3019 => to_slv(opcode_type, 16#80#),
      3020 => to_slv(opcode_type, 16#07#),
      3021 => to_slv(opcode_type, 16#05#),
      3022 => to_slv(opcode_type, 16#0D#),
      3023 => to_slv(opcode_type, 16#06#),
      3024 => to_slv(opcode_type, 16#0D#),
      3025 => to_slv(opcode_type, 16#0B#),
      3026 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#08#),
      3041 => to_slv(opcode_type, 16#01#),
      3042 => to_slv(opcode_type, 16#02#),
      3043 => to_slv(opcode_type, 16#09#),
      3044 => to_slv(opcode_type, 16#90#),
      3045 => to_slv(opcode_type, 16#0B#),
      3046 => to_slv(opcode_type, 16#06#),
      3047 => to_slv(opcode_type, 16#09#),
      3048 => to_slv(opcode_type, 16#06#),
      3049 => to_slv(opcode_type, 16#0F#),
      3050 => to_slv(opcode_type, 16#0A#),
      3051 => to_slv(opcode_type, 16#01#),
      3052 => to_slv(opcode_type, 16#10#),
      3053 => to_slv(opcode_type, 16#06#),
      3054 => to_slv(opcode_type, 16#05#),
      3055 => to_slv(opcode_type, 16#0A#),
      3056 => to_slv(opcode_type, 16#03#),
      3057 => to_slv(opcode_type, 16#0D#),
      3058 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#09#),
      3073 => to_slv(opcode_type, 16#09#),
      3074 => to_slv(opcode_type, 16#04#),
      3075 => to_slv(opcode_type, 16#02#),
      3076 => to_slv(opcode_type, 16#11#),
      3077 => to_slv(opcode_type, 16#06#),
      3078 => to_slv(opcode_type, 16#04#),
      3079 => to_slv(opcode_type, 16#37#),
      3080 => to_slv(opcode_type, 16#04#),
      3081 => to_slv(opcode_type, 16#0E#),
      3082 => to_slv(opcode_type, 16#04#),
      3083 => to_slv(opcode_type, 16#08#),
      3084 => to_slv(opcode_type, 16#08#),
      3085 => to_slv(opcode_type, 16#0F#),
      3086 => to_slv(opcode_type, 16#11#),
      3087 => to_slv(opcode_type, 16#07#),
      3088 => to_slv(opcode_type, 16#0F#),
      3089 => to_slv(opcode_type, 16#0F#),
      3090 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#06#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#03#),
      3107 => to_slv(opcode_type, 16#09#),
      3108 => to_slv(opcode_type, 16#0A#),
      3109 => to_slv(opcode_type, 16#D3#),
      3110 => to_slv(opcode_type, 16#06#),
      3111 => to_slv(opcode_type, 16#04#),
      3112 => to_slv(opcode_type, 16#0D#),
      3113 => to_slv(opcode_type, 16#03#),
      3114 => to_slv(opcode_type, 16#DF#),
      3115 => to_slv(opcode_type, 16#05#),
      3116 => to_slv(opcode_type, 16#06#),
      3117 => to_slv(opcode_type, 16#03#),
      3118 => to_slv(opcode_type, 16#0D#),
      3119 => to_slv(opcode_type, 16#07#),
      3120 => to_slv(opcode_type, 16#0E#),
      3121 => to_slv(opcode_type, 16#0B#),
      3122 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#07#),
      3137 => to_slv(opcode_type, 16#03#),
      3138 => to_slv(opcode_type, 16#02#),
      3139 => to_slv(opcode_type, 16#05#),
      3140 => to_slv(opcode_type, 16#0B#),
      3141 => to_slv(opcode_type, 16#09#),
      3142 => to_slv(opcode_type, 16#09#),
      3143 => to_slv(opcode_type, 16#05#),
      3144 => to_slv(opcode_type, 16#0B#),
      3145 => to_slv(opcode_type, 16#03#),
      3146 => to_slv(opcode_type, 16#0E#),
      3147 => to_slv(opcode_type, 16#08#),
      3148 => to_slv(opcode_type, 16#08#),
      3149 => to_slv(opcode_type, 16#0E#),
      3150 => to_slv(opcode_type, 16#0B#),
      3151 => to_slv(opcode_type, 16#09#),
      3152 => to_slv(opcode_type, 16#4A#),
      3153 => to_slv(opcode_type, 16#0C#),
      3154 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#09#),
      3169 => to_slv(opcode_type, 16#02#),
      3170 => to_slv(opcode_type, 16#01#),
      3171 => to_slv(opcode_type, 16#04#),
      3172 => to_slv(opcode_type, 16#0E#),
      3173 => to_slv(opcode_type, 16#06#),
      3174 => to_slv(opcode_type, 16#08#),
      3175 => to_slv(opcode_type, 16#07#),
      3176 => to_slv(opcode_type, 16#0D#),
      3177 => to_slv(opcode_type, 16#0F#),
      3178 => to_slv(opcode_type, 16#03#),
      3179 => to_slv(opcode_type, 16#11#),
      3180 => to_slv(opcode_type, 16#06#),
      3181 => to_slv(opcode_type, 16#09#),
      3182 => to_slv(opcode_type, 16#11#),
      3183 => to_slv(opcode_type, 16#58#),
      3184 => to_slv(opcode_type, 16#02#),
      3185 => to_slv(opcode_type, 16#0E#),
      3186 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#07#),
      3201 => to_slv(opcode_type, 16#01#),
      3202 => to_slv(opcode_type, 16#05#),
      3203 => to_slv(opcode_type, 16#05#),
      3204 => to_slv(opcode_type, 16#0B#),
      3205 => to_slv(opcode_type, 16#06#),
      3206 => to_slv(opcode_type, 16#07#),
      3207 => to_slv(opcode_type, 16#03#),
      3208 => to_slv(opcode_type, 16#E2#),
      3209 => to_slv(opcode_type, 16#02#),
      3210 => to_slv(opcode_type, 16#0F#),
      3211 => to_slv(opcode_type, 16#07#),
      3212 => to_slv(opcode_type, 16#09#),
      3213 => to_slv(opcode_type, 16#11#),
      3214 => to_slv(opcode_type, 16#11#),
      3215 => to_slv(opcode_type, 16#09#),
      3216 => to_slv(opcode_type, 16#10#),
      3217 => to_slv(opcode_type, 16#0E#),
      3218 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#05#),
      3234 => to_slv(opcode_type, 16#01#),
      3235 => to_slv(opcode_type, 16#04#),
      3236 => to_slv(opcode_type, 16#0E#),
      3237 => to_slv(opcode_type, 16#07#),
      3238 => to_slv(opcode_type, 16#09#),
      3239 => to_slv(opcode_type, 16#01#),
      3240 => to_slv(opcode_type, 16#0C#),
      3241 => to_slv(opcode_type, 16#08#),
      3242 => to_slv(opcode_type, 16#0B#),
      3243 => to_slv(opcode_type, 16#0A#),
      3244 => to_slv(opcode_type, 16#09#),
      3245 => to_slv(opcode_type, 16#07#),
      3246 => to_slv(opcode_type, 16#0C#),
      3247 => to_slv(opcode_type, 16#0C#),
      3248 => to_slv(opcode_type, 16#02#),
      3249 => to_slv(opcode_type, 16#10#),
      3250 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#08#),
      3265 => to_slv(opcode_type, 16#09#),
      3266 => to_slv(opcode_type, 16#03#),
      3267 => to_slv(opcode_type, 16#09#),
      3268 => to_slv(opcode_type, 16#0D#),
      3269 => to_slv(opcode_type, 16#0A#),
      3270 => to_slv(opcode_type, 16#08#),
      3271 => to_slv(opcode_type, 16#07#),
      3272 => to_slv(opcode_type, 16#0C#),
      3273 => to_slv(opcode_type, 16#0B#),
      3274 => to_slv(opcode_type, 16#03#),
      3275 => to_slv(opcode_type, 16#0D#),
      3276 => to_slv(opcode_type, 16#01#),
      3277 => to_slv(opcode_type, 16#07#),
      3278 => to_slv(opcode_type, 16#01#),
      3279 => to_slv(opcode_type, 16#10#),
      3280 => to_slv(opcode_type, 16#02#),
      3281 => to_slv(opcode_type, 16#10#),
      3282 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#06#),
      3297 => to_slv(opcode_type, 16#01#),
      3298 => to_slv(opcode_type, 16#08#),
      3299 => to_slv(opcode_type, 16#08#),
      3300 => to_slv(opcode_type, 16#0F#),
      3301 => to_slv(opcode_type, 16#11#),
      3302 => to_slv(opcode_type, 16#01#),
      3303 => to_slv(opcode_type, 16#0F#),
      3304 => to_slv(opcode_type, 16#08#),
      3305 => to_slv(opcode_type, 16#06#),
      3306 => to_slv(opcode_type, 16#07#),
      3307 => to_slv(opcode_type, 16#0F#),
      3308 => to_slv(opcode_type, 16#0B#),
      3309 => to_slv(opcode_type, 16#05#),
      3310 => to_slv(opcode_type, 16#11#),
      3311 => to_slv(opcode_type, 16#07#),
      3312 => to_slv(opcode_type, 16#0A#),
      3313 => to_slv(opcode_type, 16#0A#),
      3314 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#06#),
      3329 => to_slv(opcode_type, 16#07#),
      3330 => to_slv(opcode_type, 16#08#),
      3331 => to_slv(opcode_type, 16#04#),
      3332 => to_slv(opcode_type, 16#0D#),
      3333 => to_slv(opcode_type, 16#03#),
      3334 => to_slv(opcode_type, 16#10#),
      3335 => to_slv(opcode_type, 16#07#),
      3336 => to_slv(opcode_type, 16#03#),
      3337 => to_slv(opcode_type, 16#0D#),
      3338 => to_slv(opcode_type, 16#03#),
      3339 => to_slv(opcode_type, 16#0D#),
      3340 => to_slv(opcode_type, 16#05#),
      3341 => to_slv(opcode_type, 16#07#),
      3342 => to_slv(opcode_type, 16#02#),
      3343 => to_slv(opcode_type, 16#0F#),
      3344 => to_slv(opcode_type, 16#04#),
      3345 => to_slv(opcode_type, 16#0F#),
      3346 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#08#),
      3361 => to_slv(opcode_type, 16#03#),
      3362 => to_slv(opcode_type, 16#02#),
      3363 => to_slv(opcode_type, 16#06#),
      3364 => to_slv(opcode_type, 16#10#),
      3365 => to_slv(opcode_type, 16#0E#),
      3366 => to_slv(opcode_type, 16#08#),
      3367 => to_slv(opcode_type, 16#02#),
      3368 => to_slv(opcode_type, 16#07#),
      3369 => to_slv(opcode_type, 16#0F#),
      3370 => to_slv(opcode_type, 16#0E#),
      3371 => to_slv(opcode_type, 16#07#),
      3372 => to_slv(opcode_type, 16#09#),
      3373 => to_slv(opcode_type, 16#0E#),
      3374 => to_slv(opcode_type, 16#0B#),
      3375 => to_slv(opcode_type, 16#07#),
      3376 => to_slv(opcode_type, 16#0D#),
      3377 => to_slv(opcode_type, 16#10#),
      3378 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#06#),
      3393 => to_slv(opcode_type, 16#08#),
      3394 => to_slv(opcode_type, 16#03#),
      3395 => to_slv(opcode_type, 16#03#),
      3396 => to_slv(opcode_type, 16#11#),
      3397 => to_slv(opcode_type, 16#01#),
      3398 => to_slv(opcode_type, 16#04#),
      3399 => to_slv(opcode_type, 16#0A#),
      3400 => to_slv(opcode_type, 16#07#),
      3401 => to_slv(opcode_type, 16#05#),
      3402 => to_slv(opcode_type, 16#06#),
      3403 => to_slv(opcode_type, 16#11#),
      3404 => to_slv(opcode_type, 16#0F#),
      3405 => to_slv(opcode_type, 16#09#),
      3406 => to_slv(opcode_type, 16#02#),
      3407 => to_slv(opcode_type, 16#0D#),
      3408 => to_slv(opcode_type, 16#05#),
      3409 => to_slv(opcode_type, 16#0D#),
      3410 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#07#),
      3426 => to_slv(opcode_type, 16#03#),
      3427 => to_slv(opcode_type, 16#08#),
      3428 => to_slv(opcode_type, 16#0E#),
      3429 => to_slv(opcode_type, 16#0F#),
      3430 => to_slv(opcode_type, 16#04#),
      3431 => to_slv(opcode_type, 16#09#),
      3432 => to_slv(opcode_type, 16#0A#),
      3433 => to_slv(opcode_type, 16#0E#),
      3434 => to_slv(opcode_type, 16#05#),
      3435 => to_slv(opcode_type, 16#06#),
      3436 => to_slv(opcode_type, 16#08#),
      3437 => to_slv(opcode_type, 16#0E#),
      3438 => to_slv(opcode_type, 16#0E#),
      3439 => to_slv(opcode_type, 16#07#),
      3440 => to_slv(opcode_type, 16#0B#),
      3441 => to_slv(opcode_type, 16#16#),
      3442 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#08#),
      3457 => to_slv(opcode_type, 16#09#),
      3458 => to_slv(opcode_type, 16#09#),
      3459 => to_slv(opcode_type, 16#01#),
      3460 => to_slv(opcode_type, 16#0E#),
      3461 => to_slv(opcode_type, 16#05#),
      3462 => to_slv(opcode_type, 16#0D#),
      3463 => to_slv(opcode_type, 16#04#),
      3464 => to_slv(opcode_type, 16#03#),
      3465 => to_slv(opcode_type, 16#0F#),
      3466 => to_slv(opcode_type, 16#08#),
      3467 => to_slv(opcode_type, 16#03#),
      3468 => to_slv(opcode_type, 16#01#),
      3469 => to_slv(opcode_type, 16#0B#),
      3470 => to_slv(opcode_type, 16#08#),
      3471 => to_slv(opcode_type, 16#05#),
      3472 => to_slv(opcode_type, 16#0E#),
      3473 => to_slv(opcode_type, 16#53#),
      3474 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#06#),
      3489 => to_slv(opcode_type, 16#04#),
      3490 => to_slv(opcode_type, 16#03#),
      3491 => to_slv(opcode_type, 16#08#),
      3492 => to_slv(opcode_type, 16#0B#),
      3493 => to_slv(opcode_type, 16#0F#),
      3494 => to_slv(opcode_type, 16#06#),
      3495 => to_slv(opcode_type, 16#01#),
      3496 => to_slv(opcode_type, 16#09#),
      3497 => to_slv(opcode_type, 16#0D#),
      3498 => to_slv(opcode_type, 16#11#),
      3499 => to_slv(opcode_type, 16#07#),
      3500 => to_slv(opcode_type, 16#09#),
      3501 => to_slv(opcode_type, 16#0B#),
      3502 => to_slv(opcode_type, 16#11#),
      3503 => to_slv(opcode_type, 16#06#),
      3504 => to_slv(opcode_type, 16#0C#),
      3505 => to_slv(opcode_type, 16#0D#),
      3506 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#08#),
      3521 => to_slv(opcode_type, 16#02#),
      3522 => to_slv(opcode_type, 16#09#),
      3523 => to_slv(opcode_type, 16#06#),
      3524 => to_slv(opcode_type, 16#17#),
      3525 => to_slv(opcode_type, 16#10#),
      3526 => to_slv(opcode_type, 16#08#),
      3527 => to_slv(opcode_type, 16#0D#),
      3528 => to_slv(opcode_type, 16#0A#),
      3529 => to_slv(opcode_type, 16#08#),
      3530 => to_slv(opcode_type, 16#01#),
      3531 => to_slv(opcode_type, 16#08#),
      3532 => to_slv(opcode_type, 16#0C#),
      3533 => to_slv(opcode_type, 16#0D#),
      3534 => to_slv(opcode_type, 16#06#),
      3535 => to_slv(opcode_type, 16#04#),
      3536 => to_slv(opcode_type, 16#0E#),
      3537 => to_slv(opcode_type, 16#11#),
      3538 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#07#),
      3553 => to_slv(opcode_type, 16#08#),
      3554 => to_slv(opcode_type, 16#04#),
      3555 => to_slv(opcode_type, 16#07#),
      3556 => to_slv(opcode_type, 16#10#),
      3557 => to_slv(opcode_type, 16#0C#),
      3558 => to_slv(opcode_type, 16#03#),
      3559 => to_slv(opcode_type, 16#05#),
      3560 => to_slv(opcode_type, 16#0F#),
      3561 => to_slv(opcode_type, 16#08#),
      3562 => to_slv(opcode_type, 16#04#),
      3563 => to_slv(opcode_type, 16#06#),
      3564 => to_slv(opcode_type, 16#11#),
      3565 => to_slv(opcode_type, 16#23#),
      3566 => to_slv(opcode_type, 16#08#),
      3567 => to_slv(opcode_type, 16#05#),
      3568 => to_slv(opcode_type, 16#10#),
      3569 => to_slv(opcode_type, 16#10#),
      3570 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#07#),
      3585 => to_slv(opcode_type, 16#03#),
      3586 => to_slv(opcode_type, 16#06#),
      3587 => to_slv(opcode_type, 16#06#),
      3588 => to_slv(opcode_type, 16#0B#),
      3589 => to_slv(opcode_type, 16#0C#),
      3590 => to_slv(opcode_type, 16#04#),
      3591 => to_slv(opcode_type, 16#0E#),
      3592 => to_slv(opcode_type, 16#06#),
      3593 => to_slv(opcode_type, 16#07#),
      3594 => to_slv(opcode_type, 16#05#),
      3595 => to_slv(opcode_type, 16#10#),
      3596 => to_slv(opcode_type, 16#04#),
      3597 => to_slv(opcode_type, 16#0D#),
      3598 => to_slv(opcode_type, 16#08#),
      3599 => to_slv(opcode_type, 16#02#),
      3600 => to_slv(opcode_type, 16#0D#),
      3601 => to_slv(opcode_type, 16#0F#),
      3602 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#09#),
      3617 => to_slv(opcode_type, 16#09#),
      3618 => to_slv(opcode_type, 16#08#),
      3619 => to_slv(opcode_type, 16#01#),
      3620 => to_slv(opcode_type, 16#A9#),
      3621 => to_slv(opcode_type, 16#06#),
      3622 => to_slv(opcode_type, 16#90#),
      3623 => to_slv(opcode_type, 16#10#),
      3624 => to_slv(opcode_type, 16#05#),
      3625 => to_slv(opcode_type, 16#08#),
      3626 => to_slv(opcode_type, 16#10#),
      3627 => to_slv(opcode_type, 16#0D#),
      3628 => to_slv(opcode_type, 16#01#),
      3629 => to_slv(opcode_type, 16#08#),
      3630 => to_slv(opcode_type, 16#03#),
      3631 => to_slv(opcode_type, 16#0A#),
      3632 => to_slv(opcode_type, 16#03#),
      3633 => to_slv(opcode_type, 16#0D#),
      3634 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#09#),
      3649 => to_slv(opcode_type, 16#04#),
      3650 => to_slv(opcode_type, 16#05#),
      3651 => to_slv(opcode_type, 16#03#),
      3652 => to_slv(opcode_type, 16#0E#),
      3653 => to_slv(opcode_type, 16#07#),
      3654 => to_slv(opcode_type, 16#09#),
      3655 => to_slv(opcode_type, 16#06#),
      3656 => to_slv(opcode_type, 16#0C#),
      3657 => to_slv(opcode_type, 16#0E#),
      3658 => to_slv(opcode_type, 16#01#),
      3659 => to_slv(opcode_type, 16#0C#),
      3660 => to_slv(opcode_type, 16#07#),
      3661 => to_slv(opcode_type, 16#03#),
      3662 => to_slv(opcode_type, 16#0B#),
      3663 => to_slv(opcode_type, 16#08#),
      3664 => to_slv(opcode_type, 16#0C#),
      3665 => to_slv(opcode_type, 16#48#),
      3666 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#08#),
      3681 => to_slv(opcode_type, 16#01#),
      3682 => to_slv(opcode_type, 16#05#),
      3683 => to_slv(opcode_type, 16#06#),
      3684 => to_slv(opcode_type, 16#11#),
      3685 => to_slv(opcode_type, 16#10#),
      3686 => to_slv(opcode_type, 16#08#),
      3687 => to_slv(opcode_type, 16#04#),
      3688 => to_slv(opcode_type, 16#08#),
      3689 => to_slv(opcode_type, 16#0D#),
      3690 => to_slv(opcode_type, 16#0A#),
      3691 => to_slv(opcode_type, 16#08#),
      3692 => to_slv(opcode_type, 16#06#),
      3693 => to_slv(opcode_type, 16#11#),
      3694 => to_slv(opcode_type, 16#42#),
      3695 => to_slv(opcode_type, 16#09#),
      3696 => to_slv(opcode_type, 16#0B#),
      3697 => to_slv(opcode_type, 16#0F#),
      3698 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#08#),
      3713 => to_slv(opcode_type, 16#04#),
      3714 => to_slv(opcode_type, 16#07#),
      3715 => to_slv(opcode_type, 16#02#),
      3716 => to_slv(opcode_type, 16#0D#),
      3717 => to_slv(opcode_type, 16#09#),
      3718 => to_slv(opcode_type, 16#10#),
      3719 => to_slv(opcode_type, 16#0A#),
      3720 => to_slv(opcode_type, 16#07#),
      3721 => to_slv(opcode_type, 16#02#),
      3722 => to_slv(opcode_type, 16#09#),
      3723 => to_slv(opcode_type, 16#11#),
      3724 => to_slv(opcode_type, 16#0A#),
      3725 => to_slv(opcode_type, 16#06#),
      3726 => to_slv(opcode_type, 16#03#),
      3727 => to_slv(opcode_type, 16#0D#),
      3728 => to_slv(opcode_type, 16#01#),
      3729 => to_slv(opcode_type, 16#0D#),
      3730 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#07#),
      3745 => to_slv(opcode_type, 16#05#),
      3746 => to_slv(opcode_type, 16#05#),
      3747 => to_slv(opcode_type, 16#05#),
      3748 => to_slv(opcode_type, 16#10#),
      3749 => to_slv(opcode_type, 16#06#),
      3750 => to_slv(opcode_type, 16#09#),
      3751 => to_slv(opcode_type, 16#01#),
      3752 => to_slv(opcode_type, 16#0A#),
      3753 => to_slv(opcode_type, 16#08#),
      3754 => to_slv(opcode_type, 16#0D#),
      3755 => to_slv(opcode_type, 16#11#),
      3756 => to_slv(opcode_type, 16#06#),
      3757 => to_slv(opcode_type, 16#07#),
      3758 => to_slv(opcode_type, 16#0E#),
      3759 => to_slv(opcode_type, 16#0B#),
      3760 => to_slv(opcode_type, 16#01#),
      3761 => to_slv(opcode_type, 16#0D#),
      3762 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#07#),
      3777 => to_slv(opcode_type, 16#03#),
      3778 => to_slv(opcode_type, 16#03#),
      3779 => to_slv(opcode_type, 16#08#),
      3780 => to_slv(opcode_type, 16#0C#),
      3781 => to_slv(opcode_type, 16#0F#),
      3782 => to_slv(opcode_type, 16#06#),
      3783 => to_slv(opcode_type, 16#02#),
      3784 => to_slv(opcode_type, 16#06#),
      3785 => to_slv(opcode_type, 16#CA#),
      3786 => to_slv(opcode_type, 16#11#),
      3787 => to_slv(opcode_type, 16#07#),
      3788 => to_slv(opcode_type, 16#08#),
      3789 => to_slv(opcode_type, 16#0F#),
      3790 => to_slv(opcode_type, 16#0E#),
      3791 => to_slv(opcode_type, 16#09#),
      3792 => to_slv(opcode_type, 16#0B#),
      3793 => to_slv(opcode_type, 16#0F#),
      3794 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#06#),
      3809 => to_slv(opcode_type, 16#05#),
      3810 => to_slv(opcode_type, 16#06#),
      3811 => to_slv(opcode_type, 16#01#),
      3812 => to_slv(opcode_type, 16#10#),
      3813 => to_slv(opcode_type, 16#02#),
      3814 => to_slv(opcode_type, 16#0C#),
      3815 => to_slv(opcode_type, 16#06#),
      3816 => to_slv(opcode_type, 16#06#),
      3817 => to_slv(opcode_type, 16#09#),
      3818 => to_slv(opcode_type, 16#0B#),
      3819 => to_slv(opcode_type, 16#0F#),
      3820 => to_slv(opcode_type, 16#08#),
      3821 => to_slv(opcode_type, 16#10#),
      3822 => to_slv(opcode_type, 16#0B#),
      3823 => to_slv(opcode_type, 16#08#),
      3824 => to_slv(opcode_type, 16#C4#),
      3825 => to_slv(opcode_type, 16#11#),
      3826 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#08#),
      3841 => to_slv(opcode_type, 16#08#),
      3842 => to_slv(opcode_type, 16#08#),
      3843 => to_slv(opcode_type, 16#01#),
      3844 => to_slv(opcode_type, 16#10#),
      3845 => to_slv(opcode_type, 16#05#),
      3846 => to_slv(opcode_type, 16#0F#),
      3847 => to_slv(opcode_type, 16#06#),
      3848 => to_slv(opcode_type, 16#01#),
      3849 => to_slv(opcode_type, 16#0D#),
      3850 => to_slv(opcode_type, 16#02#),
      3851 => to_slv(opcode_type, 16#0E#),
      3852 => to_slv(opcode_type, 16#09#),
      3853 => to_slv(opcode_type, 16#08#),
      3854 => to_slv(opcode_type, 16#03#),
      3855 => to_slv(opcode_type, 16#0C#),
      3856 => to_slv(opcode_type, 16#0A#),
      3857 => to_slv(opcode_type, 16#11#),
      3858 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#09#),
      3873 => to_slv(opcode_type, 16#07#),
      3874 => to_slv(opcode_type, 16#03#),
      3875 => to_slv(opcode_type, 16#08#),
      3876 => to_slv(opcode_type, 16#0A#),
      3877 => to_slv(opcode_type, 16#0C#),
      3878 => to_slv(opcode_type, 16#04#),
      3879 => to_slv(opcode_type, 16#02#),
      3880 => to_slv(opcode_type, 16#0A#),
      3881 => to_slv(opcode_type, 16#08#),
      3882 => to_slv(opcode_type, 16#07#),
      3883 => to_slv(opcode_type, 16#01#),
      3884 => to_slv(opcode_type, 16#0E#),
      3885 => to_slv(opcode_type, 16#02#),
      3886 => to_slv(opcode_type, 16#10#),
      3887 => to_slv(opcode_type, 16#04#),
      3888 => to_slv(opcode_type, 16#04#),
      3889 => to_slv(opcode_type, 16#0E#),
      3890 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#07#),
      3905 => to_slv(opcode_type, 16#07#),
      3906 => to_slv(opcode_type, 16#07#),
      3907 => to_slv(opcode_type, 16#04#),
      3908 => to_slv(opcode_type, 16#0F#),
      3909 => to_slv(opcode_type, 16#09#),
      3910 => to_slv(opcode_type, 16#0B#),
      3911 => to_slv(opcode_type, 16#0F#),
      3912 => to_slv(opcode_type, 16#01#),
      3913 => to_slv(opcode_type, 16#02#),
      3914 => to_slv(opcode_type, 16#0E#),
      3915 => to_slv(opcode_type, 16#07#),
      3916 => to_slv(opcode_type, 16#08#),
      3917 => to_slv(opcode_type, 16#03#),
      3918 => to_slv(opcode_type, 16#0E#),
      3919 => to_slv(opcode_type, 16#01#),
      3920 => to_slv(opcode_type, 16#77#),
      3921 => to_slv(opcode_type, 16#0D#),
      3922 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#06#),
      3937 => to_slv(opcode_type, 16#05#),
      3938 => to_slv(opcode_type, 16#02#),
      3939 => to_slv(opcode_type, 16#03#),
      3940 => to_slv(opcode_type, 16#0D#),
      3941 => to_slv(opcode_type, 16#07#),
      3942 => to_slv(opcode_type, 16#07#),
      3943 => to_slv(opcode_type, 16#05#),
      3944 => to_slv(opcode_type, 16#0B#),
      3945 => to_slv(opcode_type, 16#07#),
      3946 => to_slv(opcode_type, 16#0F#),
      3947 => to_slv(opcode_type, 16#11#),
      3948 => to_slv(opcode_type, 16#09#),
      3949 => to_slv(opcode_type, 16#04#),
      3950 => to_slv(opcode_type, 16#0F#),
      3951 => to_slv(opcode_type, 16#09#),
      3952 => to_slv(opcode_type, 16#0A#),
      3953 => to_slv(opcode_type, 16#0F#),
      3954 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#07#),
      3969 => to_slv(opcode_type, 16#09#),
      3970 => to_slv(opcode_type, 16#08#),
      3971 => to_slv(opcode_type, 16#06#),
      3972 => to_slv(opcode_type, 16#0C#),
      3973 => to_slv(opcode_type, 16#0C#),
      3974 => to_slv(opcode_type, 16#09#),
      3975 => to_slv(opcode_type, 16#0A#),
      3976 => to_slv(opcode_type, 16#0A#),
      3977 => to_slv(opcode_type, 16#06#),
      3978 => to_slv(opcode_type, 16#05#),
      3979 => to_slv(opcode_type, 16#0A#),
      3980 => to_slv(opcode_type, 16#07#),
      3981 => to_slv(opcode_type, 16#0F#),
      3982 => to_slv(opcode_type, 16#0C#),
      3983 => to_slv(opcode_type, 16#08#),
      3984 => to_slv(opcode_type, 16#0C#),
      3985 => to_slv(opcode_type, 16#11#),
      3986 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#09#),
      4001 => to_slv(opcode_type, 16#04#),
      4002 => to_slv(opcode_type, 16#01#),
      4003 => to_slv(opcode_type, 16#02#),
      4004 => to_slv(opcode_type, 16#0A#),
      4005 => to_slv(opcode_type, 16#08#),
      4006 => to_slv(opcode_type, 16#07#),
      4007 => to_slv(opcode_type, 16#01#),
      4008 => to_slv(opcode_type, 16#11#),
      4009 => to_slv(opcode_type, 16#07#),
      4010 => to_slv(opcode_type, 16#11#),
      4011 => to_slv(opcode_type, 16#0C#),
      4012 => to_slv(opcode_type, 16#08#),
      4013 => to_slv(opcode_type, 16#06#),
      4014 => to_slv(opcode_type, 16#10#),
      4015 => to_slv(opcode_type, 16#0A#),
      4016 => to_slv(opcode_type, 16#01#),
      4017 => to_slv(opcode_type, 16#E4#),
      4018 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#06#),
      4033 => to_slv(opcode_type, 16#02#),
      4034 => to_slv(opcode_type, 16#07#),
      4035 => to_slv(opcode_type, 16#01#),
      4036 => to_slv(opcode_type, 16#0F#),
      4037 => to_slv(opcode_type, 16#06#),
      4038 => to_slv(opcode_type, 16#15#),
      4039 => to_slv(opcode_type, 16#0B#),
      4040 => to_slv(opcode_type, 16#08#),
      4041 => to_slv(opcode_type, 16#02#),
      4042 => to_slv(opcode_type, 16#05#),
      4043 => to_slv(opcode_type, 16#0D#),
      4044 => to_slv(opcode_type, 16#08#),
      4045 => to_slv(opcode_type, 16#06#),
      4046 => to_slv(opcode_type, 16#0E#),
      4047 => to_slv(opcode_type, 16#0E#),
      4048 => to_slv(opcode_type, 16#03#),
      4049 => to_slv(opcode_type, 16#0E#),
      4050 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#03#),
      4066 => to_slv(opcode_type, 16#07#),
      4067 => to_slv(opcode_type, 16#08#),
      4068 => to_slv(opcode_type, 16#DA#),
      4069 => to_slv(opcode_type, 16#11#),
      4070 => to_slv(opcode_type, 16#09#),
      4071 => to_slv(opcode_type, 16#0F#),
      4072 => to_slv(opcode_type, 16#11#),
      4073 => to_slv(opcode_type, 16#08#),
      4074 => to_slv(opcode_type, 16#02#),
      4075 => to_slv(opcode_type, 16#04#),
      4076 => to_slv(opcode_type, 16#0D#),
      4077 => to_slv(opcode_type, 16#07#),
      4078 => to_slv(opcode_type, 16#03#),
      4079 => to_slv(opcode_type, 16#0A#),
      4080 => to_slv(opcode_type, 16#02#),
      4081 => to_slv(opcode_type, 16#22#),
      4082 to 4095 => (others => '0')
  ),

    -- Bin `19`...
    18 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#06#),
      1 => to_slv(opcode_type, 16#01#),
      2 => to_slv(opcode_type, 16#07#),
      3 => to_slv(opcode_type, 16#04#),
      4 => to_slv(opcode_type, 16#0E#),
      5 => to_slv(opcode_type, 16#02#),
      6 => to_slv(opcode_type, 16#0D#),
      7 => to_slv(opcode_type, 16#09#),
      8 => to_slv(opcode_type, 16#09#),
      9 => to_slv(opcode_type, 16#03#),
      10 => to_slv(opcode_type, 16#0D#),
      11 => to_slv(opcode_type, 16#06#),
      12 => to_slv(opcode_type, 16#11#),
      13 => to_slv(opcode_type, 16#0D#),
      14 => to_slv(opcode_type, 16#08#),
      15 => to_slv(opcode_type, 16#07#),
      16 => to_slv(opcode_type, 16#0D#),
      17 => to_slv(opcode_type, 16#10#),
      18 => to_slv(opcode_type, 16#0A#),
      19 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#08#),
      33 => to_slv(opcode_type, 16#03#),
      34 => to_slv(opcode_type, 16#01#),
      35 => to_slv(opcode_type, 16#06#),
      36 => to_slv(opcode_type, 16#0B#),
      37 => to_slv(opcode_type, 16#C8#),
      38 => to_slv(opcode_type, 16#08#),
      39 => to_slv(opcode_type, 16#09#),
      40 => to_slv(opcode_type, 16#09#),
      41 => to_slv(opcode_type, 16#10#),
      42 => to_slv(opcode_type, 16#0B#),
      43 => to_slv(opcode_type, 16#07#),
      44 => to_slv(opcode_type, 16#0B#),
      45 => to_slv(opcode_type, 16#0F#),
      46 => to_slv(opcode_type, 16#09#),
      47 => to_slv(opcode_type, 16#08#),
      48 => to_slv(opcode_type, 16#10#),
      49 => to_slv(opcode_type, 16#A6#),
      50 => to_slv(opcode_type, 16#FE#),
      51 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#08#),
      65 => to_slv(opcode_type, 16#06#),
      66 => to_slv(opcode_type, 16#01#),
      67 => to_slv(opcode_type, 16#01#),
      68 => to_slv(opcode_type, 16#0F#),
      69 => to_slv(opcode_type, 16#08#),
      70 => to_slv(opcode_type, 16#07#),
      71 => to_slv(opcode_type, 16#B3#),
      72 => to_slv(opcode_type, 16#10#),
      73 => to_slv(opcode_type, 16#06#),
      74 => to_slv(opcode_type, 16#0F#),
      75 => to_slv(opcode_type, 16#0E#),
      76 => to_slv(opcode_type, 16#03#),
      77 => to_slv(opcode_type, 16#07#),
      78 => to_slv(opcode_type, 16#07#),
      79 => to_slv(opcode_type, 16#11#),
      80 => to_slv(opcode_type, 16#0F#),
      81 => to_slv(opcode_type, 16#03#),
      82 => to_slv(opcode_type, 16#0B#),
      83 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#06#),
      97 => to_slv(opcode_type, 16#04#),
      98 => to_slv(opcode_type, 16#07#),
      99 => to_slv(opcode_type, 16#02#),
      100 => to_slv(opcode_type, 16#0C#),
      101 => to_slv(opcode_type, 16#06#),
      102 => to_slv(opcode_type, 16#C0#),
      103 => to_slv(opcode_type, 16#11#),
      104 => to_slv(opcode_type, 16#09#),
      105 => to_slv(opcode_type, 16#04#),
      106 => to_slv(opcode_type, 16#05#),
      107 => to_slv(opcode_type, 16#0C#),
      108 => to_slv(opcode_type, 16#06#),
      109 => to_slv(opcode_type, 16#09#),
      110 => to_slv(opcode_type, 16#C9#),
      111 => to_slv(opcode_type, 16#0E#),
      112 => to_slv(opcode_type, 16#08#),
      113 => to_slv(opcode_type, 16#0D#),
      114 => to_slv(opcode_type, 16#11#),
      115 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#08#),
      129 => to_slv(opcode_type, 16#06#),
      130 => to_slv(opcode_type, 16#09#),
      131 => to_slv(opcode_type, 16#04#),
      132 => to_slv(opcode_type, 16#11#),
      133 => to_slv(opcode_type, 16#01#),
      134 => to_slv(opcode_type, 16#0B#),
      135 => to_slv(opcode_type, 16#09#),
      136 => to_slv(opcode_type, 16#02#),
      137 => to_slv(opcode_type, 16#10#),
      138 => to_slv(opcode_type, 16#08#),
      139 => to_slv(opcode_type, 16#10#),
      140 => to_slv(opcode_type, 16#10#),
      141 => to_slv(opcode_type, 16#01#),
      142 => to_slv(opcode_type, 16#09#),
      143 => to_slv(opcode_type, 16#02#),
      144 => to_slv(opcode_type, 16#0F#),
      145 => to_slv(opcode_type, 16#01#),
      146 => to_slv(opcode_type, 16#0A#),
      147 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#08#),
      161 => to_slv(opcode_type, 16#06#),
      162 => to_slv(opcode_type, 16#06#),
      163 => to_slv(opcode_type, 16#08#),
      164 => to_slv(opcode_type, 16#0B#),
      165 => to_slv(opcode_type, 16#0E#),
      166 => to_slv(opcode_type, 16#05#),
      167 => to_slv(opcode_type, 16#0B#),
      168 => to_slv(opcode_type, 16#06#),
      169 => to_slv(opcode_type, 16#05#),
      170 => to_slv(opcode_type, 16#C6#),
      171 => to_slv(opcode_type, 16#07#),
      172 => to_slv(opcode_type, 16#92#),
      173 => to_slv(opcode_type, 16#11#),
      174 => to_slv(opcode_type, 16#08#),
      175 => to_slv(opcode_type, 16#01#),
      176 => to_slv(opcode_type, 16#05#),
      177 => to_slv(opcode_type, 16#0D#),
      178 => to_slv(opcode_type, 16#10#),
      179 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#09#),
      193 => to_slv(opcode_type, 16#04#),
      194 => to_slv(opcode_type, 16#08#),
      195 => to_slv(opcode_type, 16#04#),
      196 => to_slv(opcode_type, 16#0F#),
      197 => to_slv(opcode_type, 16#08#),
      198 => to_slv(opcode_type, 16#11#),
      199 => to_slv(opcode_type, 16#0E#),
      200 => to_slv(opcode_type, 16#07#),
      201 => to_slv(opcode_type, 16#01#),
      202 => to_slv(opcode_type, 16#03#),
      203 => to_slv(opcode_type, 16#10#),
      204 => to_slv(opcode_type, 16#06#),
      205 => to_slv(opcode_type, 16#08#),
      206 => to_slv(opcode_type, 16#0D#),
      207 => to_slv(opcode_type, 16#0E#),
      208 => to_slv(opcode_type, 16#09#),
      209 => to_slv(opcode_type, 16#0C#),
      210 => to_slv(opcode_type, 16#0E#),
      211 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#08#),
      225 => to_slv(opcode_type, 16#02#),
      226 => to_slv(opcode_type, 16#06#),
      227 => to_slv(opcode_type, 16#09#),
      228 => to_slv(opcode_type, 16#0D#),
      229 => to_slv(opcode_type, 16#0F#),
      230 => to_slv(opcode_type, 16#07#),
      231 => to_slv(opcode_type, 16#0A#),
      232 => to_slv(opcode_type, 16#11#),
      233 => to_slv(opcode_type, 16#06#),
      234 => to_slv(opcode_type, 16#07#),
      235 => to_slv(opcode_type, 16#02#),
      236 => to_slv(opcode_type, 16#0D#),
      237 => to_slv(opcode_type, 16#07#),
      238 => to_slv(opcode_type, 16#0A#),
      239 => to_slv(opcode_type, 16#0F#),
      240 => to_slv(opcode_type, 16#08#),
      241 => to_slv(opcode_type, 16#0C#),
      242 => to_slv(opcode_type, 16#0E#),
      243 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#06#),
      257 => to_slv(opcode_type, 16#07#),
      258 => to_slv(opcode_type, 16#05#),
      259 => to_slv(opcode_type, 16#02#),
      260 => to_slv(opcode_type, 16#10#),
      261 => to_slv(opcode_type, 16#06#),
      262 => to_slv(opcode_type, 16#06#),
      263 => to_slv(opcode_type, 16#0F#),
      264 => to_slv(opcode_type, 16#0B#),
      265 => to_slv(opcode_type, 16#08#),
      266 => to_slv(opcode_type, 16#0A#),
      267 => to_slv(opcode_type, 16#0D#),
      268 => to_slv(opcode_type, 16#04#),
      269 => to_slv(opcode_type, 16#08#),
      270 => to_slv(opcode_type, 16#08#),
      271 => to_slv(opcode_type, 16#0F#),
      272 => to_slv(opcode_type, 16#10#),
      273 => to_slv(opcode_type, 16#05#),
      274 => to_slv(opcode_type, 16#A7#),
      275 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#08#),
      289 => to_slv(opcode_type, 16#07#),
      290 => to_slv(opcode_type, 16#03#),
      291 => to_slv(opcode_type, 16#05#),
      292 => to_slv(opcode_type, 16#0D#),
      293 => to_slv(opcode_type, 16#02#),
      294 => to_slv(opcode_type, 16#03#),
      295 => to_slv(opcode_type, 16#10#),
      296 => to_slv(opcode_type, 16#07#),
      297 => to_slv(opcode_type, 16#01#),
      298 => to_slv(opcode_type, 16#01#),
      299 => to_slv(opcode_type, 16#0B#),
      300 => to_slv(opcode_type, 16#07#),
      301 => to_slv(opcode_type, 16#06#),
      302 => to_slv(opcode_type, 16#10#),
      303 => to_slv(opcode_type, 16#0F#),
      304 => to_slv(opcode_type, 16#07#),
      305 => to_slv(opcode_type, 16#0C#),
      306 => to_slv(opcode_type, 16#11#),
      307 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#06#),
      321 => to_slv(opcode_type, 16#04#),
      322 => to_slv(opcode_type, 16#05#),
      323 => to_slv(opcode_type, 16#06#),
      324 => to_slv(opcode_type, 16#D9#),
      325 => to_slv(opcode_type, 16#F3#),
      326 => to_slv(opcode_type, 16#07#),
      327 => to_slv(opcode_type, 16#07#),
      328 => to_slv(opcode_type, 16#06#),
      329 => to_slv(opcode_type, 16#11#),
      330 => to_slv(opcode_type, 16#0C#),
      331 => to_slv(opcode_type, 16#04#),
      332 => to_slv(opcode_type, 16#0F#),
      333 => to_slv(opcode_type, 16#09#),
      334 => to_slv(opcode_type, 16#08#),
      335 => to_slv(opcode_type, 16#0D#),
      336 => to_slv(opcode_type, 16#0A#),
      337 => to_slv(opcode_type, 16#05#),
      338 => to_slv(opcode_type, 16#0C#),
      339 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#06#),
      353 => to_slv(opcode_type, 16#09#),
      354 => to_slv(opcode_type, 16#09#),
      355 => to_slv(opcode_type, 16#01#),
      356 => to_slv(opcode_type, 16#0C#),
      357 => to_slv(opcode_type, 16#01#),
      358 => to_slv(opcode_type, 16#10#),
      359 => to_slv(opcode_type, 16#05#),
      360 => to_slv(opcode_type, 16#06#),
      361 => to_slv(opcode_type, 16#EC#),
      362 => to_slv(opcode_type, 16#0B#),
      363 => to_slv(opcode_type, 16#04#),
      364 => to_slv(opcode_type, 16#06#),
      365 => to_slv(opcode_type, 16#07#),
      366 => to_slv(opcode_type, 16#10#),
      367 => to_slv(opcode_type, 16#E0#),
      368 => to_slv(opcode_type, 16#08#),
      369 => to_slv(opcode_type, 16#0C#),
      370 => to_slv(opcode_type, 16#0D#),
      371 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#09#),
      385 => to_slv(opcode_type, 16#08#),
      386 => to_slv(opcode_type, 16#08#),
      387 => to_slv(opcode_type, 16#04#),
      388 => to_slv(opcode_type, 16#0D#),
      389 => to_slv(opcode_type, 16#08#),
      390 => to_slv(opcode_type, 16#11#),
      391 => to_slv(opcode_type, 16#11#),
      392 => to_slv(opcode_type, 16#09#),
      393 => to_slv(opcode_type, 16#05#),
      394 => to_slv(opcode_type, 16#0C#),
      395 => to_slv(opcode_type, 16#06#),
      396 => to_slv(opcode_type, 16#0A#),
      397 => to_slv(opcode_type, 16#0F#),
      398 => to_slv(opcode_type, 16#07#),
      399 => to_slv(opcode_type, 16#03#),
      400 => to_slv(opcode_type, 16#03#),
      401 => to_slv(opcode_type, 16#0A#),
      402 => to_slv(opcode_type, 16#10#),
      403 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#07#),
      417 => to_slv(opcode_type, 16#02#),
      418 => to_slv(opcode_type, 16#02#),
      419 => to_slv(opcode_type, 16#04#),
      420 => to_slv(opcode_type, 16#0E#),
      421 => to_slv(opcode_type, 16#06#),
      422 => to_slv(opcode_type, 16#09#),
      423 => to_slv(opcode_type, 16#07#),
      424 => to_slv(opcode_type, 16#0F#),
      425 => to_slv(opcode_type, 16#0D#),
      426 => to_slv(opcode_type, 16#06#),
      427 => to_slv(opcode_type, 16#11#),
      428 => to_slv(opcode_type, 16#0E#),
      429 => to_slv(opcode_type, 16#08#),
      430 => to_slv(opcode_type, 16#07#),
      431 => to_slv(opcode_type, 16#0A#),
      432 => to_slv(opcode_type, 16#0B#),
      433 => to_slv(opcode_type, 16#05#),
      434 => to_slv(opcode_type, 16#0C#),
      435 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#06#),
      449 => to_slv(opcode_type, 16#04#),
      450 => to_slv(opcode_type, 16#06#),
      451 => to_slv(opcode_type, 16#01#),
      452 => to_slv(opcode_type, 16#0D#),
      453 => to_slv(opcode_type, 16#03#),
      454 => to_slv(opcode_type, 16#0B#),
      455 => to_slv(opcode_type, 16#09#),
      456 => to_slv(opcode_type, 16#05#),
      457 => to_slv(opcode_type, 16#09#),
      458 => to_slv(opcode_type, 16#0B#),
      459 => to_slv(opcode_type, 16#0D#),
      460 => to_slv(opcode_type, 16#09#),
      461 => to_slv(opcode_type, 16#09#),
      462 => to_slv(opcode_type, 16#0A#),
      463 => to_slv(opcode_type, 16#0E#),
      464 => to_slv(opcode_type, 16#08#),
      465 => to_slv(opcode_type, 16#0D#),
      466 => to_slv(opcode_type, 16#72#),
      467 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#08#),
      481 => to_slv(opcode_type, 16#08#),
      482 => to_slv(opcode_type, 16#03#),
      483 => to_slv(opcode_type, 16#01#),
      484 => to_slv(opcode_type, 16#11#),
      485 => to_slv(opcode_type, 16#05#),
      486 => to_slv(opcode_type, 16#03#),
      487 => to_slv(opcode_type, 16#10#),
      488 => to_slv(opcode_type, 16#07#),
      489 => to_slv(opcode_type, 16#01#),
      490 => to_slv(opcode_type, 16#09#),
      491 => to_slv(opcode_type, 16#0B#),
      492 => to_slv(opcode_type, 16#0A#),
      493 => to_slv(opcode_type, 16#08#),
      494 => to_slv(opcode_type, 16#04#),
      495 => to_slv(opcode_type, 16#0F#),
      496 => to_slv(opcode_type, 16#06#),
      497 => to_slv(opcode_type, 16#0E#),
      498 => to_slv(opcode_type, 16#0F#),
      499 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#08#),
      513 => to_slv(opcode_type, 16#06#),
      514 => to_slv(opcode_type, 16#05#),
      515 => to_slv(opcode_type, 16#02#),
      516 => to_slv(opcode_type, 16#10#),
      517 => to_slv(opcode_type, 16#01#),
      518 => to_slv(opcode_type, 16#09#),
      519 => to_slv(opcode_type, 16#0D#),
      520 => to_slv(opcode_type, 16#0D#),
      521 => to_slv(opcode_type, 16#09#),
      522 => to_slv(opcode_type, 16#01#),
      523 => to_slv(opcode_type, 16#08#),
      524 => to_slv(opcode_type, 16#58#),
      525 => to_slv(opcode_type, 16#0A#),
      526 => to_slv(opcode_type, 16#09#),
      527 => to_slv(opcode_type, 16#01#),
      528 => to_slv(opcode_type, 16#0A#),
      529 => to_slv(opcode_type, 16#03#),
      530 => to_slv(opcode_type, 16#0B#),
      531 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#08#),
      545 => to_slv(opcode_type, 16#03#),
      546 => to_slv(opcode_type, 16#06#),
      547 => to_slv(opcode_type, 16#05#),
      548 => to_slv(opcode_type, 16#0A#),
      549 => to_slv(opcode_type, 16#02#),
      550 => to_slv(opcode_type, 16#0E#),
      551 => to_slv(opcode_type, 16#06#),
      552 => to_slv(opcode_type, 16#07#),
      553 => to_slv(opcode_type, 16#09#),
      554 => to_slv(opcode_type, 16#10#),
      555 => to_slv(opcode_type, 16#0A#),
      556 => to_slv(opcode_type, 16#09#),
      557 => to_slv(opcode_type, 16#0E#),
      558 => to_slv(opcode_type, 16#11#),
      559 => to_slv(opcode_type, 16#05#),
      560 => to_slv(opcode_type, 16#07#),
      561 => to_slv(opcode_type, 16#0A#),
      562 => to_slv(opcode_type, 16#0A#),
      563 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#06#),
      577 => to_slv(opcode_type, 16#06#),
      578 => to_slv(opcode_type, 16#04#),
      579 => to_slv(opcode_type, 16#09#),
      580 => to_slv(opcode_type, 16#0E#),
      581 => to_slv(opcode_type, 16#0F#),
      582 => to_slv(opcode_type, 16#09#),
      583 => to_slv(opcode_type, 16#01#),
      584 => to_slv(opcode_type, 16#10#),
      585 => to_slv(opcode_type, 16#09#),
      586 => to_slv(opcode_type, 16#0F#),
      587 => to_slv(opcode_type, 16#37#),
      588 => to_slv(opcode_type, 16#08#),
      589 => to_slv(opcode_type, 16#06#),
      590 => to_slv(opcode_type, 16#09#),
      591 => to_slv(opcode_type, 16#10#),
      592 => to_slv(opcode_type, 16#0D#),
      593 => to_slv(opcode_type, 16#0C#),
      594 => to_slv(opcode_type, 16#10#),
      595 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#06#),
      609 => to_slv(opcode_type, 16#08#),
      610 => to_slv(opcode_type, 16#09#),
      611 => to_slv(opcode_type, 16#06#),
      612 => to_slv(opcode_type, 16#0A#),
      613 => to_slv(opcode_type, 16#0D#),
      614 => to_slv(opcode_type, 16#07#),
      615 => to_slv(opcode_type, 16#0F#),
      616 => to_slv(opcode_type, 16#0C#),
      617 => to_slv(opcode_type, 16#04#),
      618 => to_slv(opcode_type, 16#04#),
      619 => to_slv(opcode_type, 16#0E#),
      620 => to_slv(opcode_type, 16#06#),
      621 => to_slv(opcode_type, 16#04#),
      622 => to_slv(opcode_type, 16#05#),
      623 => to_slv(opcode_type, 16#10#),
      624 => to_slv(opcode_type, 16#05#),
      625 => to_slv(opcode_type, 16#04#),
      626 => to_slv(opcode_type, 16#0D#),
      627 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#09#),
      641 => to_slv(opcode_type, 16#02#),
      642 => to_slv(opcode_type, 16#02#),
      643 => to_slv(opcode_type, 16#09#),
      644 => to_slv(opcode_type, 16#0B#),
      645 => to_slv(opcode_type, 16#0B#),
      646 => to_slv(opcode_type, 16#08#),
      647 => to_slv(opcode_type, 16#09#),
      648 => to_slv(opcode_type, 16#01#),
      649 => to_slv(opcode_type, 16#48#),
      650 => to_slv(opcode_type, 16#08#),
      651 => to_slv(opcode_type, 16#0B#),
      652 => to_slv(opcode_type, 16#11#),
      653 => to_slv(opcode_type, 16#06#),
      654 => to_slv(opcode_type, 16#08#),
      655 => to_slv(opcode_type, 16#11#),
      656 => to_slv(opcode_type, 16#11#),
      657 => to_slv(opcode_type, 16#03#),
      658 => to_slv(opcode_type, 16#0D#),
      659 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#06#),
      673 => to_slv(opcode_type, 16#01#),
      674 => to_slv(opcode_type, 16#05#),
      675 => to_slv(opcode_type, 16#08#),
      676 => to_slv(opcode_type, 16#0B#),
      677 => to_slv(opcode_type, 16#0C#),
      678 => to_slv(opcode_type, 16#06#),
      679 => to_slv(opcode_type, 16#06#),
      680 => to_slv(opcode_type, 16#04#),
      681 => to_slv(opcode_type, 16#10#),
      682 => to_slv(opcode_type, 16#06#),
      683 => to_slv(opcode_type, 16#0D#),
      684 => to_slv(opcode_type, 16#0B#),
      685 => to_slv(opcode_type, 16#09#),
      686 => to_slv(opcode_type, 16#09#),
      687 => to_slv(opcode_type, 16#0E#),
      688 => to_slv(opcode_type, 16#0C#),
      689 => to_slv(opcode_type, 16#04#),
      690 => to_slv(opcode_type, 16#0F#),
      691 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#09#),
      705 => to_slv(opcode_type, 16#08#),
      706 => to_slv(opcode_type, 16#04#),
      707 => to_slv(opcode_type, 16#01#),
      708 => to_slv(opcode_type, 16#10#),
      709 => to_slv(opcode_type, 16#09#),
      710 => to_slv(opcode_type, 16#09#),
      711 => to_slv(opcode_type, 16#0A#),
      712 => to_slv(opcode_type, 16#0A#),
      713 => to_slv(opcode_type, 16#07#),
      714 => to_slv(opcode_type, 16#0F#),
      715 => to_slv(opcode_type, 16#0B#),
      716 => to_slv(opcode_type, 16#03#),
      717 => to_slv(opcode_type, 16#06#),
      718 => to_slv(opcode_type, 16#05#),
      719 => to_slv(opcode_type, 16#0F#),
      720 => to_slv(opcode_type, 16#09#),
      721 => to_slv(opcode_type, 16#0A#),
      722 => to_slv(opcode_type, 16#0D#),
      723 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#09#),
      737 => to_slv(opcode_type, 16#05#),
      738 => to_slv(opcode_type, 16#09#),
      739 => to_slv(opcode_type, 16#03#),
      740 => to_slv(opcode_type, 16#0C#),
      741 => to_slv(opcode_type, 16#06#),
      742 => to_slv(opcode_type, 16#0E#),
      743 => to_slv(opcode_type, 16#0E#),
      744 => to_slv(opcode_type, 16#06#),
      745 => to_slv(opcode_type, 16#06#),
      746 => to_slv(opcode_type, 16#08#),
      747 => to_slv(opcode_type, 16#0D#),
      748 => to_slv(opcode_type, 16#0A#),
      749 => to_slv(opcode_type, 16#02#),
      750 => to_slv(opcode_type, 16#10#),
      751 => to_slv(opcode_type, 16#08#),
      752 => to_slv(opcode_type, 16#02#),
      753 => to_slv(opcode_type, 16#0F#),
      754 => to_slv(opcode_type, 16#0F#),
      755 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#06#),
      769 => to_slv(opcode_type, 16#02#),
      770 => to_slv(opcode_type, 16#04#),
      771 => to_slv(opcode_type, 16#07#),
      772 => to_slv(opcode_type, 16#E0#),
      773 => to_slv(opcode_type, 16#0B#),
      774 => to_slv(opcode_type, 16#09#),
      775 => to_slv(opcode_type, 16#07#),
      776 => to_slv(opcode_type, 16#07#),
      777 => to_slv(opcode_type, 16#10#),
      778 => to_slv(opcode_type, 16#0A#),
      779 => to_slv(opcode_type, 16#08#),
      780 => to_slv(opcode_type, 16#10#),
      781 => to_slv(opcode_type, 16#0A#),
      782 => to_slv(opcode_type, 16#09#),
      783 => to_slv(opcode_type, 16#04#),
      784 => to_slv(opcode_type, 16#0B#),
      785 => to_slv(opcode_type, 16#04#),
      786 => to_slv(opcode_type, 16#0F#),
      787 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#09#),
      801 => to_slv(opcode_type, 16#05#),
      802 => to_slv(opcode_type, 16#08#),
      803 => to_slv(opcode_type, 16#01#),
      804 => to_slv(opcode_type, 16#0C#),
      805 => to_slv(opcode_type, 16#07#),
      806 => to_slv(opcode_type, 16#0B#),
      807 => to_slv(opcode_type, 16#0B#),
      808 => to_slv(opcode_type, 16#09#),
      809 => to_slv(opcode_type, 16#04#),
      810 => to_slv(opcode_type, 16#08#),
      811 => to_slv(opcode_type, 16#0E#),
      812 => to_slv(opcode_type, 16#10#),
      813 => to_slv(opcode_type, 16#08#),
      814 => to_slv(opcode_type, 16#08#),
      815 => to_slv(opcode_type, 16#11#),
      816 => to_slv(opcode_type, 16#0C#),
      817 => to_slv(opcode_type, 16#01#),
      818 => to_slv(opcode_type, 16#0B#),
      819 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#07#),
      833 => to_slv(opcode_type, 16#04#),
      834 => to_slv(opcode_type, 16#02#),
      835 => to_slv(opcode_type, 16#09#),
      836 => to_slv(opcode_type, 16#FA#),
      837 => to_slv(opcode_type, 16#0C#),
      838 => to_slv(opcode_type, 16#07#),
      839 => to_slv(opcode_type, 16#07#),
      840 => to_slv(opcode_type, 16#04#),
      841 => to_slv(opcode_type, 16#10#),
      842 => to_slv(opcode_type, 16#04#),
      843 => to_slv(opcode_type, 16#0D#),
      844 => to_slv(opcode_type, 16#07#),
      845 => to_slv(opcode_type, 16#06#),
      846 => to_slv(opcode_type, 16#0E#),
      847 => to_slv(opcode_type, 16#0F#),
      848 => to_slv(opcode_type, 16#08#),
      849 => to_slv(opcode_type, 16#7B#),
      850 => to_slv(opcode_type, 16#10#),
      851 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#07#),
      865 => to_slv(opcode_type, 16#05#),
      866 => to_slv(opcode_type, 16#02#),
      867 => to_slv(opcode_type, 16#07#),
      868 => to_slv(opcode_type, 16#0F#),
      869 => to_slv(opcode_type, 16#0E#),
      870 => to_slv(opcode_type, 16#07#),
      871 => to_slv(opcode_type, 16#07#),
      872 => to_slv(opcode_type, 16#08#),
      873 => to_slv(opcode_type, 16#0B#),
      874 => to_slv(opcode_type, 16#11#),
      875 => to_slv(opcode_type, 16#09#),
      876 => to_slv(opcode_type, 16#11#),
      877 => to_slv(opcode_type, 16#10#),
      878 => to_slv(opcode_type, 16#07#),
      879 => to_slv(opcode_type, 16#01#),
      880 => to_slv(opcode_type, 16#0D#),
      881 => to_slv(opcode_type, 16#02#),
      882 => to_slv(opcode_type, 16#0F#),
      883 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#01#),
      898 => to_slv(opcode_type, 16#09#),
      899 => to_slv(opcode_type, 16#06#),
      900 => to_slv(opcode_type, 16#0D#),
      901 => to_slv(opcode_type, 16#6B#),
      902 => to_slv(opcode_type, 16#06#),
      903 => to_slv(opcode_type, 16#0E#),
      904 => to_slv(opcode_type, 16#0C#),
      905 => to_slv(opcode_type, 16#08#),
      906 => to_slv(opcode_type, 16#07#),
      907 => to_slv(opcode_type, 16#08#),
      908 => to_slv(opcode_type, 16#10#),
      909 => to_slv(opcode_type, 16#10#),
      910 => to_slv(opcode_type, 16#03#),
      911 => to_slv(opcode_type, 16#1E#),
      912 => to_slv(opcode_type, 16#01#),
      913 => to_slv(opcode_type, 16#04#),
      914 => to_slv(opcode_type, 16#0A#),
      915 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#08#),
      929 => to_slv(opcode_type, 16#08#),
      930 => to_slv(opcode_type, 16#09#),
      931 => to_slv(opcode_type, 16#09#),
      932 => to_slv(opcode_type, 16#0B#),
      933 => to_slv(opcode_type, 16#10#),
      934 => to_slv(opcode_type, 16#08#),
      935 => to_slv(opcode_type, 16#0A#),
      936 => to_slv(opcode_type, 16#0F#),
      937 => to_slv(opcode_type, 16#08#),
      938 => to_slv(opcode_type, 16#08#),
      939 => to_slv(opcode_type, 16#49#),
      940 => to_slv(opcode_type, 16#11#),
      941 => to_slv(opcode_type, 16#05#),
      942 => to_slv(opcode_type, 16#0B#),
      943 => to_slv(opcode_type, 16#09#),
      944 => to_slv(opcode_type, 16#03#),
      945 => to_slv(opcode_type, 16#10#),
      946 => to_slv(opcode_type, 16#0B#),
      947 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#03#),
      962 => to_slv(opcode_type, 16#09#),
      963 => to_slv(opcode_type, 16#01#),
      964 => to_slv(opcode_type, 16#11#),
      965 => to_slv(opcode_type, 16#09#),
      966 => to_slv(opcode_type, 16#0B#),
      967 => to_slv(opcode_type, 16#63#),
      968 => to_slv(opcode_type, 16#07#),
      969 => to_slv(opcode_type, 16#06#),
      970 => to_slv(opcode_type, 16#03#),
      971 => to_slv(opcode_type, 16#0B#),
      972 => to_slv(opcode_type, 16#03#),
      973 => to_slv(opcode_type, 16#0B#),
      974 => to_slv(opcode_type, 16#06#),
      975 => to_slv(opcode_type, 16#08#),
      976 => to_slv(opcode_type, 16#0E#),
      977 => to_slv(opcode_type, 16#0F#),
      978 => to_slv(opcode_type, 16#10#),
      979 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#09#),
      993 => to_slv(opcode_type, 16#05#),
      994 => to_slv(opcode_type, 16#07#),
      995 => to_slv(opcode_type, 16#07#),
      996 => to_slv(opcode_type, 16#0F#),
      997 => to_slv(opcode_type, 16#10#),
      998 => to_slv(opcode_type, 16#05#),
      999 => to_slv(opcode_type, 16#F3#),
      1000 => to_slv(opcode_type, 16#09#),
      1001 => to_slv(opcode_type, 16#05#),
      1002 => to_slv(opcode_type, 16#09#),
      1003 => to_slv(opcode_type, 16#11#),
      1004 => to_slv(opcode_type, 16#0A#),
      1005 => to_slv(opcode_type, 16#06#),
      1006 => to_slv(opcode_type, 16#04#),
      1007 => to_slv(opcode_type, 16#0D#),
      1008 => to_slv(opcode_type, 16#06#),
      1009 => to_slv(opcode_type, 16#10#),
      1010 => to_slv(opcode_type, 16#FC#),
      1011 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#06#),
      1025 => to_slv(opcode_type, 16#01#),
      1026 => to_slv(opcode_type, 16#04#),
      1027 => to_slv(opcode_type, 16#08#),
      1028 => to_slv(opcode_type, 16#0E#),
      1029 => to_slv(opcode_type, 16#11#),
      1030 => to_slv(opcode_type, 16#06#),
      1031 => to_slv(opcode_type, 16#07#),
      1032 => to_slv(opcode_type, 16#03#),
      1033 => to_slv(opcode_type, 16#0D#),
      1034 => to_slv(opcode_type, 16#04#),
      1035 => to_slv(opcode_type, 16#0E#),
      1036 => to_slv(opcode_type, 16#06#),
      1037 => to_slv(opcode_type, 16#08#),
      1038 => to_slv(opcode_type, 16#0D#),
      1039 => to_slv(opcode_type, 16#0E#),
      1040 => to_slv(opcode_type, 16#09#),
      1041 => to_slv(opcode_type, 16#0F#),
      1042 => to_slv(opcode_type, 16#11#),
      1043 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#08#),
      1057 => to_slv(opcode_type, 16#05#),
      1058 => to_slv(opcode_type, 16#09#),
      1059 => to_slv(opcode_type, 16#03#),
      1060 => to_slv(opcode_type, 16#0B#),
      1061 => to_slv(opcode_type, 16#07#),
      1062 => to_slv(opcode_type, 16#0C#),
      1063 => to_slv(opcode_type, 16#85#),
      1064 => to_slv(opcode_type, 16#08#),
      1065 => to_slv(opcode_type, 16#05#),
      1066 => to_slv(opcode_type, 16#07#),
      1067 => to_slv(opcode_type, 16#10#),
      1068 => to_slv(opcode_type, 16#11#),
      1069 => to_slv(opcode_type, 16#08#),
      1070 => to_slv(opcode_type, 16#05#),
      1071 => to_slv(opcode_type, 16#0C#),
      1072 => to_slv(opcode_type, 16#06#),
      1073 => to_slv(opcode_type, 16#0E#),
      1074 => to_slv(opcode_type, 16#0F#),
      1075 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#07#),
      1089 => to_slv(opcode_type, 16#05#),
      1090 => to_slv(opcode_type, 16#07#),
      1091 => to_slv(opcode_type, 16#01#),
      1092 => to_slv(opcode_type, 16#11#),
      1093 => to_slv(opcode_type, 16#04#),
      1094 => to_slv(opcode_type, 16#0D#),
      1095 => to_slv(opcode_type, 16#08#),
      1096 => to_slv(opcode_type, 16#08#),
      1097 => to_slv(opcode_type, 16#02#),
      1098 => to_slv(opcode_type, 16#0B#),
      1099 => to_slv(opcode_type, 16#05#),
      1100 => to_slv(opcode_type, 16#0C#),
      1101 => to_slv(opcode_type, 16#08#),
      1102 => to_slv(opcode_type, 16#09#),
      1103 => to_slv(opcode_type, 16#0F#),
      1104 => to_slv(opcode_type, 16#0E#),
      1105 => to_slv(opcode_type, 16#01#),
      1106 => to_slv(opcode_type, 16#11#),
      1107 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#09#),
      1121 => to_slv(opcode_type, 16#01#),
      1122 => to_slv(opcode_type, 16#05#),
      1123 => to_slv(opcode_type, 16#09#),
      1124 => to_slv(opcode_type, 16#11#),
      1125 => to_slv(opcode_type, 16#0A#),
      1126 => to_slv(opcode_type, 16#08#),
      1127 => to_slv(opcode_type, 16#06#),
      1128 => to_slv(opcode_type, 16#06#),
      1129 => to_slv(opcode_type, 16#11#),
      1130 => to_slv(opcode_type, 16#0D#),
      1131 => to_slv(opcode_type, 16#02#),
      1132 => to_slv(opcode_type, 16#0C#),
      1133 => to_slv(opcode_type, 16#07#),
      1134 => to_slv(opcode_type, 16#03#),
      1135 => to_slv(opcode_type, 16#0A#),
      1136 => to_slv(opcode_type, 16#08#),
      1137 => to_slv(opcode_type, 16#11#),
      1138 => to_slv(opcode_type, 16#0B#),
      1139 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#07#),
      1153 => to_slv(opcode_type, 16#01#),
      1154 => to_slv(opcode_type, 16#05#),
      1155 => to_slv(opcode_type, 16#06#),
      1156 => to_slv(opcode_type, 16#0B#),
      1157 => to_slv(opcode_type, 16#10#),
      1158 => to_slv(opcode_type, 16#09#),
      1159 => to_slv(opcode_type, 16#08#),
      1160 => to_slv(opcode_type, 16#04#),
      1161 => to_slv(opcode_type, 16#0A#),
      1162 => to_slv(opcode_type, 16#02#),
      1163 => to_slv(opcode_type, 16#0C#),
      1164 => to_slv(opcode_type, 16#06#),
      1165 => to_slv(opcode_type, 16#09#),
      1166 => to_slv(opcode_type, 16#0B#),
      1167 => to_slv(opcode_type, 16#0D#),
      1168 => to_slv(opcode_type, 16#09#),
      1169 => to_slv(opcode_type, 16#10#),
      1170 => to_slv(opcode_type, 16#0A#),
      1171 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#07#),
      1185 => to_slv(opcode_type, 16#04#),
      1186 => to_slv(opcode_type, 16#03#),
      1187 => to_slv(opcode_type, 16#04#),
      1188 => to_slv(opcode_type, 16#0F#),
      1189 => to_slv(opcode_type, 16#09#),
      1190 => to_slv(opcode_type, 16#07#),
      1191 => to_slv(opcode_type, 16#02#),
      1192 => to_slv(opcode_type, 16#0D#),
      1193 => to_slv(opcode_type, 16#09#),
      1194 => to_slv(opcode_type, 16#0F#),
      1195 => to_slv(opcode_type, 16#0E#),
      1196 => to_slv(opcode_type, 16#07#),
      1197 => to_slv(opcode_type, 16#08#),
      1198 => to_slv(opcode_type, 16#10#),
      1199 => to_slv(opcode_type, 16#0F#),
      1200 => to_slv(opcode_type, 16#06#),
      1201 => to_slv(opcode_type, 16#0B#),
      1202 => to_slv(opcode_type, 16#0D#),
      1203 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#08#),
      1217 => to_slv(opcode_type, 16#06#),
      1218 => to_slv(opcode_type, 16#08#),
      1219 => to_slv(opcode_type, 16#08#),
      1220 => to_slv(opcode_type, 16#11#),
      1221 => to_slv(opcode_type, 16#10#),
      1222 => to_slv(opcode_type, 16#03#),
      1223 => to_slv(opcode_type, 16#10#),
      1224 => to_slv(opcode_type, 16#07#),
      1225 => to_slv(opcode_type, 16#02#),
      1226 => to_slv(opcode_type, 16#0B#),
      1227 => to_slv(opcode_type, 16#02#),
      1228 => to_slv(opcode_type, 16#0D#),
      1229 => to_slv(opcode_type, 16#08#),
      1230 => to_slv(opcode_type, 16#09#),
      1231 => to_slv(opcode_type, 16#05#),
      1232 => to_slv(opcode_type, 16#0C#),
      1233 => to_slv(opcode_type, 16#0D#),
      1234 => to_slv(opcode_type, 16#11#),
      1235 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#06#),
      1249 => to_slv(opcode_type, 16#09#),
      1250 => to_slv(opcode_type, 16#06#),
      1251 => to_slv(opcode_type, 16#06#),
      1252 => to_slv(opcode_type, 16#0B#),
      1253 => to_slv(opcode_type, 16#0E#),
      1254 => to_slv(opcode_type, 16#02#),
      1255 => to_slv(opcode_type, 16#0A#),
      1256 => to_slv(opcode_type, 16#03#),
      1257 => to_slv(opcode_type, 16#05#),
      1258 => to_slv(opcode_type, 16#11#),
      1259 => to_slv(opcode_type, 16#08#),
      1260 => to_slv(opcode_type, 16#03#),
      1261 => to_slv(opcode_type, 16#04#),
      1262 => to_slv(opcode_type, 16#0D#),
      1263 => to_slv(opcode_type, 16#09#),
      1264 => to_slv(opcode_type, 16#04#),
      1265 => to_slv(opcode_type, 16#0F#),
      1266 => to_slv(opcode_type, 16#0E#),
      1267 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#01#),
      1282 => to_slv(opcode_type, 16#01#),
      1283 => to_slv(opcode_type, 16#08#),
      1284 => to_slv(opcode_type, 16#10#),
      1285 => to_slv(opcode_type, 16#0C#),
      1286 => to_slv(opcode_type, 16#06#),
      1287 => to_slv(opcode_type, 16#09#),
      1288 => to_slv(opcode_type, 16#01#),
      1289 => to_slv(opcode_type, 16#0C#),
      1290 => to_slv(opcode_type, 16#09#),
      1291 => to_slv(opcode_type, 16#0E#),
      1292 => to_slv(opcode_type, 16#11#),
      1293 => to_slv(opcode_type, 16#07#),
      1294 => to_slv(opcode_type, 16#06#),
      1295 => to_slv(opcode_type, 16#E7#),
      1296 => to_slv(opcode_type, 16#0D#),
      1297 => to_slv(opcode_type, 16#03#),
      1298 => to_slv(opcode_type, 16#10#),
      1299 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#07#),
      1313 => to_slv(opcode_type, 16#01#),
      1314 => to_slv(opcode_type, 16#03#),
      1315 => to_slv(opcode_type, 16#04#),
      1316 => to_slv(opcode_type, 16#0C#),
      1317 => to_slv(opcode_type, 16#08#),
      1318 => to_slv(opcode_type, 16#08#),
      1319 => to_slv(opcode_type, 16#03#),
      1320 => to_slv(opcode_type, 16#10#),
      1321 => to_slv(opcode_type, 16#06#),
      1322 => to_slv(opcode_type, 16#0D#),
      1323 => to_slv(opcode_type, 16#10#),
      1324 => to_slv(opcode_type, 16#07#),
      1325 => to_slv(opcode_type, 16#06#),
      1326 => to_slv(opcode_type, 16#11#),
      1327 => to_slv(opcode_type, 16#0A#),
      1328 => to_slv(opcode_type, 16#06#),
      1329 => to_slv(opcode_type, 16#0F#),
      1330 => to_slv(opcode_type, 16#0C#),
      1331 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#09#),
      1345 => to_slv(opcode_type, 16#05#),
      1346 => to_slv(opcode_type, 16#04#),
      1347 => to_slv(opcode_type, 16#01#),
      1348 => to_slv(opcode_type, 16#0C#),
      1349 => to_slv(opcode_type, 16#06#),
      1350 => to_slv(opcode_type, 16#08#),
      1351 => to_slv(opcode_type, 16#06#),
      1352 => to_slv(opcode_type, 16#10#),
      1353 => to_slv(opcode_type, 16#11#),
      1354 => to_slv(opcode_type, 16#09#),
      1355 => to_slv(opcode_type, 16#FD#),
      1356 => to_slv(opcode_type, 16#0E#),
      1357 => to_slv(opcode_type, 16#07#),
      1358 => to_slv(opcode_type, 16#04#),
      1359 => to_slv(opcode_type, 16#0F#),
      1360 => to_slv(opcode_type, 16#08#),
      1361 => to_slv(opcode_type, 16#10#),
      1362 => to_slv(opcode_type, 16#11#),
      1363 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#07#),
      1377 => to_slv(opcode_type, 16#09#),
      1378 => to_slv(opcode_type, 16#07#),
      1379 => to_slv(opcode_type, 16#08#),
      1380 => to_slv(opcode_type, 16#0C#),
      1381 => to_slv(opcode_type, 16#10#),
      1382 => to_slv(opcode_type, 16#01#),
      1383 => to_slv(opcode_type, 16#0F#),
      1384 => to_slv(opcode_type, 16#01#),
      1385 => to_slv(opcode_type, 16#04#),
      1386 => to_slv(opcode_type, 16#10#),
      1387 => to_slv(opcode_type, 16#01#),
      1388 => to_slv(opcode_type, 16#08#),
      1389 => to_slv(opcode_type, 16#08#),
      1390 => to_slv(opcode_type, 16#0C#),
      1391 => to_slv(opcode_type, 16#0D#),
      1392 => to_slv(opcode_type, 16#08#),
      1393 => to_slv(opcode_type, 16#0A#),
      1394 => to_slv(opcode_type, 16#0A#),
      1395 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#06#),
      1410 => to_slv(opcode_type, 16#09#),
      1411 => to_slv(opcode_type, 16#01#),
      1412 => to_slv(opcode_type, 16#0A#),
      1413 => to_slv(opcode_type, 16#02#),
      1414 => to_slv(opcode_type, 16#0D#),
      1415 => to_slv(opcode_type, 16#02#),
      1416 => to_slv(opcode_type, 16#01#),
      1417 => to_slv(opcode_type, 16#0D#),
      1418 => to_slv(opcode_type, 16#06#),
      1419 => to_slv(opcode_type, 16#08#),
      1420 => to_slv(opcode_type, 16#05#),
      1421 => to_slv(opcode_type, 16#0B#),
      1422 => to_slv(opcode_type, 16#02#),
      1423 => to_slv(opcode_type, 16#10#),
      1424 => to_slv(opcode_type, 16#01#),
      1425 => to_slv(opcode_type, 16#03#),
      1426 => to_slv(opcode_type, 16#0E#),
      1427 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#09#),
      1441 => to_slv(opcode_type, 16#07#),
      1442 => to_slv(opcode_type, 16#03#),
      1443 => to_slv(opcode_type, 16#09#),
      1444 => to_slv(opcode_type, 16#0E#),
      1445 => to_slv(opcode_type, 16#0A#),
      1446 => to_slv(opcode_type, 16#09#),
      1447 => to_slv(opcode_type, 16#01#),
      1448 => to_slv(opcode_type, 16#0F#),
      1449 => to_slv(opcode_type, 16#01#),
      1450 => to_slv(opcode_type, 16#0C#),
      1451 => to_slv(opcode_type, 16#05#),
      1452 => to_slv(opcode_type, 16#09#),
      1453 => to_slv(opcode_type, 16#09#),
      1454 => to_slv(opcode_type, 16#0F#),
      1455 => to_slv(opcode_type, 16#8F#),
      1456 => to_slv(opcode_type, 16#07#),
      1457 => to_slv(opcode_type, 16#0D#),
      1458 => to_slv(opcode_type, 16#11#),
      1459 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#07#),
      1473 => to_slv(opcode_type, 16#04#),
      1474 => to_slv(opcode_type, 16#08#),
      1475 => to_slv(opcode_type, 16#02#),
      1476 => to_slv(opcode_type, 16#11#),
      1477 => to_slv(opcode_type, 16#08#),
      1478 => to_slv(opcode_type, 16#10#),
      1479 => to_slv(opcode_type, 16#0E#),
      1480 => to_slv(opcode_type, 16#07#),
      1481 => to_slv(opcode_type, 16#03#),
      1482 => to_slv(opcode_type, 16#09#),
      1483 => to_slv(opcode_type, 16#11#),
      1484 => to_slv(opcode_type, 16#11#),
      1485 => to_slv(opcode_type, 16#06#),
      1486 => to_slv(opcode_type, 16#06#),
      1487 => to_slv(opcode_type, 16#0B#),
      1488 => to_slv(opcode_type, 16#10#),
      1489 => to_slv(opcode_type, 16#03#),
      1490 => to_slv(opcode_type, 16#0F#),
      1491 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#06#),
      1505 => to_slv(opcode_type, 16#08#),
      1506 => to_slv(opcode_type, 16#08#),
      1507 => to_slv(opcode_type, 16#09#),
      1508 => to_slv(opcode_type, 16#11#),
      1509 => to_slv(opcode_type, 16#0F#),
      1510 => to_slv(opcode_type, 16#03#),
      1511 => to_slv(opcode_type, 16#0D#),
      1512 => to_slv(opcode_type, 16#02#),
      1513 => to_slv(opcode_type, 16#04#),
      1514 => to_slv(opcode_type, 16#0E#),
      1515 => to_slv(opcode_type, 16#02#),
      1516 => to_slv(opcode_type, 16#09#),
      1517 => to_slv(opcode_type, 16#06#),
      1518 => to_slv(opcode_type, 16#0C#),
      1519 => to_slv(opcode_type, 16#E5#),
      1520 => to_slv(opcode_type, 16#09#),
      1521 => to_slv(opcode_type, 16#2C#),
      1522 => to_slv(opcode_type, 16#0A#),
      1523 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#06#),
      1537 => to_slv(opcode_type, 16#02#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#05#),
      1540 => to_slv(opcode_type, 16#0E#),
      1541 => to_slv(opcode_type, 16#06#),
      1542 => to_slv(opcode_type, 16#10#),
      1543 => to_slv(opcode_type, 16#0E#),
      1544 => to_slv(opcode_type, 16#08#),
      1545 => to_slv(opcode_type, 16#07#),
      1546 => to_slv(opcode_type, 16#03#),
      1547 => to_slv(opcode_type, 16#10#),
      1548 => to_slv(opcode_type, 16#01#),
      1549 => to_slv(opcode_type, 16#0F#),
      1550 => to_slv(opcode_type, 16#08#),
      1551 => to_slv(opcode_type, 16#04#),
      1552 => to_slv(opcode_type, 16#0D#),
      1553 => to_slv(opcode_type, 16#03#),
      1554 => to_slv(opcode_type, 16#0F#),
      1555 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#07#),
      1569 => to_slv(opcode_type, 16#05#),
      1570 => to_slv(opcode_type, 16#06#),
      1571 => to_slv(opcode_type, 16#08#),
      1572 => to_slv(opcode_type, 16#0E#),
      1573 => to_slv(opcode_type, 16#0A#),
      1574 => to_slv(opcode_type, 16#09#),
      1575 => to_slv(opcode_type, 16#0F#),
      1576 => to_slv(opcode_type, 16#0D#),
      1577 => to_slv(opcode_type, 16#06#),
      1578 => to_slv(opcode_type, 16#03#),
      1579 => to_slv(opcode_type, 16#05#),
      1580 => to_slv(opcode_type, 16#0B#),
      1581 => to_slv(opcode_type, 16#06#),
      1582 => to_slv(opcode_type, 16#02#),
      1583 => to_slv(opcode_type, 16#0C#),
      1584 => to_slv(opcode_type, 16#09#),
      1585 => to_slv(opcode_type, 16#0E#),
      1586 => to_slv(opcode_type, 16#0D#),
      1587 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#03#),
      1602 => to_slv(opcode_type, 16#06#),
      1603 => to_slv(opcode_type, 16#07#),
      1604 => to_slv(opcode_type, 16#11#),
      1605 => to_slv(opcode_type, 16#0A#),
      1606 => to_slv(opcode_type, 16#09#),
      1607 => to_slv(opcode_type, 16#0E#),
      1608 => to_slv(opcode_type, 16#0E#),
      1609 => to_slv(opcode_type, 16#07#),
      1610 => to_slv(opcode_type, 16#04#),
      1611 => to_slv(opcode_type, 16#01#),
      1612 => to_slv(opcode_type, 16#11#),
      1613 => to_slv(opcode_type, 16#06#),
      1614 => to_slv(opcode_type, 16#08#),
      1615 => to_slv(opcode_type, 16#0A#),
      1616 => to_slv(opcode_type, 16#0E#),
      1617 => to_slv(opcode_type, 16#05#),
      1618 => to_slv(opcode_type, 16#0C#),
      1619 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#07#),
      1633 => to_slv(opcode_type, 16#07#),
      1634 => to_slv(opcode_type, 16#05#),
      1635 => to_slv(opcode_type, 16#03#),
      1636 => to_slv(opcode_type, 16#0D#),
      1637 => to_slv(opcode_type, 16#07#),
      1638 => to_slv(opcode_type, 16#01#),
      1639 => to_slv(opcode_type, 16#0D#),
      1640 => to_slv(opcode_type, 16#09#),
      1641 => to_slv(opcode_type, 16#11#),
      1642 => to_slv(opcode_type, 16#0D#),
      1643 => to_slv(opcode_type, 16#02#),
      1644 => to_slv(opcode_type, 16#07#),
      1645 => to_slv(opcode_type, 16#08#),
      1646 => to_slv(opcode_type, 16#0C#),
      1647 => to_slv(opcode_type, 16#0A#),
      1648 => to_slv(opcode_type, 16#07#),
      1649 => to_slv(opcode_type, 16#0A#),
      1650 => to_slv(opcode_type, 16#0C#),
      1651 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#06#),
      1665 => to_slv(opcode_type, 16#05#),
      1666 => to_slv(opcode_type, 16#09#),
      1667 => to_slv(opcode_type, 16#02#),
      1668 => to_slv(opcode_type, 16#0E#),
      1669 => to_slv(opcode_type, 16#03#),
      1670 => to_slv(opcode_type, 16#10#),
      1671 => to_slv(opcode_type, 16#08#),
      1672 => to_slv(opcode_type, 16#08#),
      1673 => to_slv(opcode_type, 16#07#),
      1674 => to_slv(opcode_type, 16#11#),
      1675 => to_slv(opcode_type, 16#11#),
      1676 => to_slv(opcode_type, 16#08#),
      1677 => to_slv(opcode_type, 16#0E#),
      1678 => to_slv(opcode_type, 16#EA#),
      1679 => to_slv(opcode_type, 16#06#),
      1680 => to_slv(opcode_type, 16#02#),
      1681 => to_slv(opcode_type, 16#0A#),
      1682 => to_slv(opcode_type, 16#0E#),
      1683 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#09#),
      1697 => to_slv(opcode_type, 16#02#),
      1698 => to_slv(opcode_type, 16#07#),
      1699 => to_slv(opcode_type, 16#03#),
      1700 => to_slv(opcode_type, 16#11#),
      1701 => to_slv(opcode_type, 16#05#),
      1702 => to_slv(opcode_type, 16#0B#),
      1703 => to_slv(opcode_type, 16#09#),
      1704 => to_slv(opcode_type, 16#05#),
      1705 => to_slv(opcode_type, 16#06#),
      1706 => to_slv(opcode_type, 16#0C#),
      1707 => to_slv(opcode_type, 16#10#),
      1708 => to_slv(opcode_type, 16#08#),
      1709 => to_slv(opcode_type, 16#09#),
      1710 => to_slv(opcode_type, 16#10#),
      1711 => to_slv(opcode_type, 16#0E#),
      1712 => to_slv(opcode_type, 16#08#),
      1713 => to_slv(opcode_type, 16#0C#),
      1714 => to_slv(opcode_type, 16#0A#),
      1715 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#08#),
      1729 => to_slv(opcode_type, 16#04#),
      1730 => to_slv(opcode_type, 16#06#),
      1731 => to_slv(opcode_type, 16#04#),
      1732 => to_slv(opcode_type, 16#0F#),
      1733 => to_slv(opcode_type, 16#04#),
      1734 => to_slv(opcode_type, 16#0D#),
      1735 => to_slv(opcode_type, 16#09#),
      1736 => to_slv(opcode_type, 16#07#),
      1737 => to_slv(opcode_type, 16#07#),
      1738 => to_slv(opcode_type, 16#FF#),
      1739 => to_slv(opcode_type, 16#0D#),
      1740 => to_slv(opcode_type, 16#09#),
      1741 => to_slv(opcode_type, 16#11#),
      1742 => to_slv(opcode_type, 16#0F#),
      1743 => to_slv(opcode_type, 16#03#),
      1744 => to_slv(opcode_type, 16#08#),
      1745 => to_slv(opcode_type, 16#10#),
      1746 => to_slv(opcode_type, 16#0F#),
      1747 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#09#),
      1761 => to_slv(opcode_type, 16#09#),
      1762 => to_slv(opcode_type, 16#03#),
      1763 => to_slv(opcode_type, 16#09#),
      1764 => to_slv(opcode_type, 16#0E#),
      1765 => to_slv(opcode_type, 16#0B#),
      1766 => to_slv(opcode_type, 16#02#),
      1767 => to_slv(opcode_type, 16#02#),
      1768 => to_slv(opcode_type, 16#10#),
      1769 => to_slv(opcode_type, 16#07#),
      1770 => to_slv(opcode_type, 16#02#),
      1771 => to_slv(opcode_type, 16#03#),
      1772 => to_slv(opcode_type, 16#10#),
      1773 => to_slv(opcode_type, 16#06#),
      1774 => to_slv(opcode_type, 16#09#),
      1775 => to_slv(opcode_type, 16#0E#),
      1776 => to_slv(opcode_type, 16#0B#),
      1777 => to_slv(opcode_type, 16#02#),
      1778 => to_slv(opcode_type, 16#10#),
      1779 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#08#),
      1793 => to_slv(opcode_type, 16#02#),
      1794 => to_slv(opcode_type, 16#06#),
      1795 => to_slv(opcode_type, 16#03#),
      1796 => to_slv(opcode_type, 16#10#),
      1797 => to_slv(opcode_type, 16#03#),
      1798 => to_slv(opcode_type, 16#0B#),
      1799 => to_slv(opcode_type, 16#06#),
      1800 => to_slv(opcode_type, 16#07#),
      1801 => to_slv(opcode_type, 16#01#),
      1802 => to_slv(opcode_type, 16#11#),
      1803 => to_slv(opcode_type, 16#06#),
      1804 => to_slv(opcode_type, 16#0E#),
      1805 => to_slv(opcode_type, 16#96#),
      1806 => to_slv(opcode_type, 16#09#),
      1807 => to_slv(opcode_type, 16#05#),
      1808 => to_slv(opcode_type, 16#0C#),
      1809 => to_slv(opcode_type, 16#04#),
      1810 => to_slv(opcode_type, 16#0A#),
      1811 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#06#),
      1825 => to_slv(opcode_type, 16#01#),
      1826 => to_slv(opcode_type, 16#07#),
      1827 => to_slv(opcode_type, 16#02#),
      1828 => to_slv(opcode_type, 16#0D#),
      1829 => to_slv(opcode_type, 16#08#),
      1830 => to_slv(opcode_type, 16#0A#),
      1831 => to_slv(opcode_type, 16#0D#),
      1832 => to_slv(opcode_type, 16#07#),
      1833 => to_slv(opcode_type, 16#06#),
      1834 => to_slv(opcode_type, 16#06#),
      1835 => to_slv(opcode_type, 16#11#),
      1836 => to_slv(opcode_type, 16#10#),
      1837 => to_slv(opcode_type, 16#02#),
      1838 => to_slv(opcode_type, 16#0C#),
      1839 => to_slv(opcode_type, 16#05#),
      1840 => to_slv(opcode_type, 16#09#),
      1841 => to_slv(opcode_type, 16#0B#),
      1842 => to_slv(opcode_type, 16#0A#),
      1843 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#06#),
      1857 => to_slv(opcode_type, 16#06#),
      1858 => to_slv(opcode_type, 16#07#),
      1859 => to_slv(opcode_type, 16#02#),
      1860 => to_slv(opcode_type, 16#0E#),
      1861 => to_slv(opcode_type, 16#07#),
      1862 => to_slv(opcode_type, 16#0E#),
      1863 => to_slv(opcode_type, 16#0B#),
      1864 => to_slv(opcode_type, 16#08#),
      1865 => to_slv(opcode_type, 16#07#),
      1866 => to_slv(opcode_type, 16#11#),
      1867 => to_slv(opcode_type, 16#0F#),
      1868 => to_slv(opcode_type, 16#01#),
      1869 => to_slv(opcode_type, 16#0D#),
      1870 => to_slv(opcode_type, 16#09#),
      1871 => to_slv(opcode_type, 16#04#),
      1872 => to_slv(opcode_type, 16#05#),
      1873 => to_slv(opcode_type, 16#10#),
      1874 => to_slv(opcode_type, 16#11#),
      1875 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#07#),
      1889 => to_slv(opcode_type, 16#05#),
      1890 => to_slv(opcode_type, 16#07#),
      1891 => to_slv(opcode_type, 16#07#),
      1892 => to_slv(opcode_type, 16#0E#),
      1893 => to_slv(opcode_type, 16#0E#),
      1894 => to_slv(opcode_type, 16#06#),
      1895 => to_slv(opcode_type, 16#10#),
      1896 => to_slv(opcode_type, 16#10#),
      1897 => to_slv(opcode_type, 16#07#),
      1898 => to_slv(opcode_type, 16#09#),
      1899 => to_slv(opcode_type, 16#05#),
      1900 => to_slv(opcode_type, 16#0B#),
      1901 => to_slv(opcode_type, 16#06#),
      1902 => to_slv(opcode_type, 16#0A#),
      1903 => to_slv(opcode_type, 16#0D#),
      1904 => to_slv(opcode_type, 16#06#),
      1905 => to_slv(opcode_type, 16#0F#),
      1906 => to_slv(opcode_type, 16#11#),
      1907 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#07#),
      1921 => to_slv(opcode_type, 16#03#),
      1922 => to_slv(opcode_type, 16#09#),
      1923 => to_slv(opcode_type, 16#09#),
      1924 => to_slv(opcode_type, 16#10#),
      1925 => to_slv(opcode_type, 16#0A#),
      1926 => to_slv(opcode_type, 16#06#),
      1927 => to_slv(opcode_type, 16#0E#),
      1928 => to_slv(opcode_type, 16#D7#),
      1929 => to_slv(opcode_type, 16#08#),
      1930 => to_slv(opcode_type, 16#07#),
      1931 => to_slv(opcode_type, 16#01#),
      1932 => to_slv(opcode_type, 16#0B#),
      1933 => to_slv(opcode_type, 16#05#),
      1934 => to_slv(opcode_type, 16#0F#),
      1935 => to_slv(opcode_type, 16#06#),
      1936 => to_slv(opcode_type, 16#05#),
      1937 => to_slv(opcode_type, 16#0C#),
      1938 => to_slv(opcode_type, 16#11#),
      1939 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#09#),
      1953 => to_slv(opcode_type, 16#03#),
      1954 => to_slv(opcode_type, 16#04#),
      1955 => to_slv(opcode_type, 16#07#),
      1956 => to_slv(opcode_type, 16#0E#),
      1957 => to_slv(opcode_type, 16#11#),
      1958 => to_slv(opcode_type, 16#06#),
      1959 => to_slv(opcode_type, 16#07#),
      1960 => to_slv(opcode_type, 16#04#),
      1961 => to_slv(opcode_type, 16#0E#),
      1962 => to_slv(opcode_type, 16#06#),
      1963 => to_slv(opcode_type, 16#0E#),
      1964 => to_slv(opcode_type, 16#0C#),
      1965 => to_slv(opcode_type, 16#07#),
      1966 => to_slv(opcode_type, 16#04#),
      1967 => to_slv(opcode_type, 16#0B#),
      1968 => to_slv(opcode_type, 16#08#),
      1969 => to_slv(opcode_type, 16#11#),
      1970 => to_slv(opcode_type, 16#0C#),
      1971 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#08#),
      1985 => to_slv(opcode_type, 16#05#),
      1986 => to_slv(opcode_type, 16#09#),
      1987 => to_slv(opcode_type, 16#07#),
      1988 => to_slv(opcode_type, 16#0E#),
      1989 => to_slv(opcode_type, 16#0C#),
      1990 => to_slv(opcode_type, 16#01#),
      1991 => to_slv(opcode_type, 16#0A#),
      1992 => to_slv(opcode_type, 16#07#),
      1993 => to_slv(opcode_type, 16#03#),
      1994 => to_slv(opcode_type, 16#04#),
      1995 => to_slv(opcode_type, 16#0B#),
      1996 => to_slv(opcode_type, 16#06#),
      1997 => to_slv(opcode_type, 16#09#),
      1998 => to_slv(opcode_type, 16#10#),
      1999 => to_slv(opcode_type, 16#0C#),
      2000 => to_slv(opcode_type, 16#09#),
      2001 => to_slv(opcode_type, 16#11#),
      2002 => to_slv(opcode_type, 16#10#),
      2003 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#09#),
      2017 => to_slv(opcode_type, 16#01#),
      2018 => to_slv(opcode_type, 16#06#),
      2019 => to_slv(opcode_type, 16#07#),
      2020 => to_slv(opcode_type, 16#0F#),
      2021 => to_slv(opcode_type, 16#0B#),
      2022 => to_slv(opcode_type, 16#05#),
      2023 => to_slv(opcode_type, 16#0C#),
      2024 => to_slv(opcode_type, 16#08#),
      2025 => to_slv(opcode_type, 16#05#),
      2026 => to_slv(opcode_type, 16#03#),
      2027 => to_slv(opcode_type, 16#0F#),
      2028 => to_slv(opcode_type, 16#06#),
      2029 => to_slv(opcode_type, 16#06#),
      2030 => to_slv(opcode_type, 16#0E#),
      2031 => to_slv(opcode_type, 16#0D#),
      2032 => to_slv(opcode_type, 16#07#),
      2033 => to_slv(opcode_type, 16#10#),
      2034 => to_slv(opcode_type, 16#0C#),
      2035 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#07#),
      2049 => to_slv(opcode_type, 16#03#),
      2050 => to_slv(opcode_type, 16#08#),
      2051 => to_slv(opcode_type, 16#03#),
      2052 => to_slv(opcode_type, 16#0F#),
      2053 => to_slv(opcode_type, 16#09#),
      2054 => to_slv(opcode_type, 16#0B#),
      2055 => to_slv(opcode_type, 16#11#),
      2056 => to_slv(opcode_type, 16#07#),
      2057 => to_slv(opcode_type, 16#08#),
      2058 => to_slv(opcode_type, 16#06#),
      2059 => to_slv(opcode_type, 16#0B#),
      2060 => to_slv(opcode_type, 16#59#),
      2061 => to_slv(opcode_type, 16#06#),
      2062 => to_slv(opcode_type, 16#11#),
      2063 => to_slv(opcode_type, 16#0E#),
      2064 => to_slv(opcode_type, 16#09#),
      2065 => to_slv(opcode_type, 16#0E#),
      2066 => to_slv(opcode_type, 16#B8#),
      2067 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#09#),
      2081 => to_slv(opcode_type, 16#02#),
      2082 => to_slv(opcode_type, 16#03#),
      2083 => to_slv(opcode_type, 16#02#),
      2084 => to_slv(opcode_type, 16#0B#),
      2085 => to_slv(opcode_type, 16#07#),
      2086 => to_slv(opcode_type, 16#06#),
      2087 => to_slv(opcode_type, 16#09#),
      2088 => to_slv(opcode_type, 16#0F#),
      2089 => to_slv(opcode_type, 16#11#),
      2090 => to_slv(opcode_type, 16#06#),
      2091 => to_slv(opcode_type, 16#0C#),
      2092 => to_slv(opcode_type, 16#11#),
      2093 => to_slv(opcode_type, 16#09#),
      2094 => to_slv(opcode_type, 16#04#),
      2095 => to_slv(opcode_type, 16#0D#),
      2096 => to_slv(opcode_type, 16#08#),
      2097 => to_slv(opcode_type, 16#0A#),
      2098 => to_slv(opcode_type, 16#0A#),
      2099 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#07#),
      2113 => to_slv(opcode_type, 16#02#),
      2114 => to_slv(opcode_type, 16#09#),
      2115 => to_slv(opcode_type, 16#07#),
      2116 => to_slv(opcode_type, 16#11#),
      2117 => to_slv(opcode_type, 16#10#),
      2118 => to_slv(opcode_type, 16#03#),
      2119 => to_slv(opcode_type, 16#0C#),
      2120 => to_slv(opcode_type, 16#09#),
      2121 => to_slv(opcode_type, 16#04#),
      2122 => to_slv(opcode_type, 16#07#),
      2123 => to_slv(opcode_type, 16#0A#),
      2124 => to_slv(opcode_type, 16#11#),
      2125 => to_slv(opcode_type, 16#08#),
      2126 => to_slv(opcode_type, 16#02#),
      2127 => to_slv(opcode_type, 16#0B#),
      2128 => to_slv(opcode_type, 16#09#),
      2129 => to_slv(opcode_type, 16#11#),
      2130 => to_slv(opcode_type, 16#0C#),
      2131 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#07#),
      2145 => to_slv(opcode_type, 16#09#),
      2146 => to_slv(opcode_type, 16#04#),
      2147 => to_slv(opcode_type, 16#02#),
      2148 => to_slv(opcode_type, 16#0B#),
      2149 => to_slv(opcode_type, 16#09#),
      2150 => to_slv(opcode_type, 16#09#),
      2151 => to_slv(opcode_type, 16#0C#),
      2152 => to_slv(opcode_type, 16#0B#),
      2153 => to_slv(opcode_type, 16#06#),
      2154 => to_slv(opcode_type, 16#0D#),
      2155 => to_slv(opcode_type, 16#0F#),
      2156 => to_slv(opcode_type, 16#01#),
      2157 => to_slv(opcode_type, 16#06#),
      2158 => to_slv(opcode_type, 16#09#),
      2159 => to_slv(opcode_type, 16#0C#),
      2160 => to_slv(opcode_type, 16#10#),
      2161 => to_slv(opcode_type, 16#05#),
      2162 => to_slv(opcode_type, 16#10#),
      2163 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#07#),
      2177 => to_slv(opcode_type, 16#06#),
      2178 => to_slv(opcode_type, 16#09#),
      2179 => to_slv(opcode_type, 16#04#),
      2180 => to_slv(opcode_type, 16#0D#),
      2181 => to_slv(opcode_type, 16#08#),
      2182 => to_slv(opcode_type, 16#0A#),
      2183 => to_slv(opcode_type, 16#0B#),
      2184 => to_slv(opcode_type, 16#01#),
      2185 => to_slv(opcode_type, 16#01#),
      2186 => to_slv(opcode_type, 16#0C#),
      2187 => to_slv(opcode_type, 16#01#),
      2188 => to_slv(opcode_type, 16#06#),
      2189 => to_slv(opcode_type, 16#07#),
      2190 => to_slv(opcode_type, 16#0A#),
      2191 => to_slv(opcode_type, 16#11#),
      2192 => to_slv(opcode_type, 16#06#),
      2193 => to_slv(opcode_type, 16#C7#),
      2194 => to_slv(opcode_type, 16#26#),
      2195 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#08#),
      2209 => to_slv(opcode_type, 16#08#),
      2210 => to_slv(opcode_type, 16#04#),
      2211 => to_slv(opcode_type, 16#05#),
      2212 => to_slv(opcode_type, 16#0C#),
      2213 => to_slv(opcode_type, 16#07#),
      2214 => to_slv(opcode_type, 16#06#),
      2215 => to_slv(opcode_type, 16#F7#),
      2216 => to_slv(opcode_type, 16#0D#),
      2217 => to_slv(opcode_type, 16#05#),
      2218 => to_slv(opcode_type, 16#0B#),
      2219 => to_slv(opcode_type, 16#07#),
      2220 => to_slv(opcode_type, 16#03#),
      2221 => to_slv(opcode_type, 16#01#),
      2222 => to_slv(opcode_type, 16#11#),
      2223 => to_slv(opcode_type, 16#01#),
      2224 => to_slv(opcode_type, 16#09#),
      2225 => to_slv(opcode_type, 16#0F#),
      2226 => to_slv(opcode_type, 16#0B#),
      2227 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#07#),
      2241 => to_slv(opcode_type, 16#04#),
      2242 => to_slv(opcode_type, 16#05#),
      2243 => to_slv(opcode_type, 16#07#),
      2244 => to_slv(opcode_type, 16#10#),
      2245 => to_slv(opcode_type, 16#10#),
      2246 => to_slv(opcode_type, 16#06#),
      2247 => to_slv(opcode_type, 16#06#),
      2248 => to_slv(opcode_type, 16#02#),
      2249 => to_slv(opcode_type, 16#0F#),
      2250 => to_slv(opcode_type, 16#07#),
      2251 => to_slv(opcode_type, 16#0B#),
      2252 => to_slv(opcode_type, 16#11#),
      2253 => to_slv(opcode_type, 16#08#),
      2254 => to_slv(opcode_type, 16#05#),
      2255 => to_slv(opcode_type, 16#0D#),
      2256 => to_slv(opcode_type, 16#07#),
      2257 => to_slv(opcode_type, 16#10#),
      2258 => to_slv(opcode_type, 16#0A#),
      2259 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#07#),
      2273 => to_slv(opcode_type, 16#03#),
      2274 => to_slv(opcode_type, 16#06#),
      2275 => to_slv(opcode_type, 16#08#),
      2276 => to_slv(opcode_type, 16#11#),
      2277 => to_slv(opcode_type, 16#0C#),
      2278 => to_slv(opcode_type, 16#03#),
      2279 => to_slv(opcode_type, 16#CB#),
      2280 => to_slv(opcode_type, 16#06#),
      2281 => to_slv(opcode_type, 16#09#),
      2282 => to_slv(opcode_type, 16#09#),
      2283 => to_slv(opcode_type, 16#0B#),
      2284 => to_slv(opcode_type, 16#0E#),
      2285 => to_slv(opcode_type, 16#06#),
      2286 => to_slv(opcode_type, 16#0B#),
      2287 => to_slv(opcode_type, 16#10#),
      2288 => to_slv(opcode_type, 16#09#),
      2289 => to_slv(opcode_type, 16#11#),
      2290 => to_slv(opcode_type, 16#10#),
      2291 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#08#),
      2305 => to_slv(opcode_type, 16#02#),
      2306 => to_slv(opcode_type, 16#07#),
      2307 => to_slv(opcode_type, 16#02#),
      2308 => to_slv(opcode_type, 16#0E#),
      2309 => to_slv(opcode_type, 16#06#),
      2310 => to_slv(opcode_type, 16#0C#),
      2311 => to_slv(opcode_type, 16#0D#),
      2312 => to_slv(opcode_type, 16#07#),
      2313 => to_slv(opcode_type, 16#09#),
      2314 => to_slv(opcode_type, 16#08#),
      2315 => to_slv(opcode_type, 16#0E#),
      2316 => to_slv(opcode_type, 16#0E#),
      2317 => to_slv(opcode_type, 16#08#),
      2318 => to_slv(opcode_type, 16#0D#),
      2319 => to_slv(opcode_type, 16#0D#),
      2320 => to_slv(opcode_type, 16#03#),
      2321 => to_slv(opcode_type, 16#03#),
      2322 => to_slv(opcode_type, 16#D5#),
      2323 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#07#),
      2337 => to_slv(opcode_type, 16#06#),
      2338 => to_slv(opcode_type, 16#04#),
      2339 => to_slv(opcode_type, 16#09#),
      2340 => to_slv(opcode_type, 16#10#),
      2341 => to_slv(opcode_type, 16#0B#),
      2342 => to_slv(opcode_type, 16#01#),
      2343 => to_slv(opcode_type, 16#02#),
      2344 => to_slv(opcode_type, 16#0C#),
      2345 => to_slv(opcode_type, 16#08#),
      2346 => to_slv(opcode_type, 16#09#),
      2347 => to_slv(opcode_type, 16#03#),
      2348 => to_slv(opcode_type, 16#0D#),
      2349 => to_slv(opcode_type, 16#02#),
      2350 => to_slv(opcode_type, 16#0B#),
      2351 => to_slv(opcode_type, 16#05#),
      2352 => to_slv(opcode_type, 16#06#),
      2353 => to_slv(opcode_type, 16#0D#),
      2354 => to_slv(opcode_type, 16#0E#),
      2355 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#09#),
      2369 => to_slv(opcode_type, 16#09#),
      2370 => to_slv(opcode_type, 16#07#),
      2371 => to_slv(opcode_type, 16#07#),
      2372 => to_slv(opcode_type, 16#B4#),
      2373 => to_slv(opcode_type, 16#0B#),
      2374 => to_slv(opcode_type, 16#05#),
      2375 => to_slv(opcode_type, 16#0B#),
      2376 => to_slv(opcode_type, 16#04#),
      2377 => to_slv(opcode_type, 16#07#),
      2378 => to_slv(opcode_type, 16#0F#),
      2379 => to_slv(opcode_type, 16#11#),
      2380 => to_slv(opcode_type, 16#09#),
      2381 => to_slv(opcode_type, 16#03#),
      2382 => to_slv(opcode_type, 16#08#),
      2383 => to_slv(opcode_type, 16#11#),
      2384 => to_slv(opcode_type, 16#0D#),
      2385 => to_slv(opcode_type, 16#05#),
      2386 => to_slv(opcode_type, 16#11#),
      2387 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#07#),
      2401 => to_slv(opcode_type, 16#09#),
      2402 => to_slv(opcode_type, 16#06#),
      2403 => to_slv(opcode_type, 16#06#),
      2404 => to_slv(opcode_type, 16#10#),
      2405 => to_slv(opcode_type, 16#0D#),
      2406 => to_slv(opcode_type, 16#02#),
      2407 => to_slv(opcode_type, 16#11#),
      2408 => to_slv(opcode_type, 16#04#),
      2409 => to_slv(opcode_type, 16#06#),
      2410 => to_slv(opcode_type, 16#4C#),
      2411 => to_slv(opcode_type, 16#0A#),
      2412 => to_slv(opcode_type, 16#05#),
      2413 => to_slv(opcode_type, 16#06#),
      2414 => to_slv(opcode_type, 16#08#),
      2415 => to_slv(opcode_type, 16#0B#),
      2416 => to_slv(opcode_type, 16#0D#),
      2417 => to_slv(opcode_type, 16#05#),
      2418 => to_slv(opcode_type, 16#10#),
      2419 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#07#),
      2433 => to_slv(opcode_type, 16#08#),
      2434 => to_slv(opcode_type, 16#04#),
      2435 => to_slv(opcode_type, 16#02#),
      2436 => to_slv(opcode_type, 16#11#),
      2437 => to_slv(opcode_type, 16#08#),
      2438 => to_slv(opcode_type, 16#03#),
      2439 => to_slv(opcode_type, 16#10#),
      2440 => to_slv(opcode_type, 16#03#),
      2441 => to_slv(opcode_type, 16#0E#),
      2442 => to_slv(opcode_type, 16#06#),
      2443 => to_slv(opcode_type, 16#07#),
      2444 => to_slv(opcode_type, 16#09#),
      2445 => to_slv(opcode_type, 16#0A#),
      2446 => to_slv(opcode_type, 16#11#),
      2447 => to_slv(opcode_type, 16#01#),
      2448 => to_slv(opcode_type, 16#CF#),
      2449 => to_slv(opcode_type, 16#02#),
      2450 => to_slv(opcode_type, 16#0D#),
      2451 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#06#),
      2465 => to_slv(opcode_type, 16#03#),
      2466 => to_slv(opcode_type, 16#01#),
      2467 => to_slv(opcode_type, 16#04#),
      2468 => to_slv(opcode_type, 16#0E#),
      2469 => to_slv(opcode_type, 16#08#),
      2470 => to_slv(opcode_type, 16#07#),
      2471 => to_slv(opcode_type, 16#03#),
      2472 => to_slv(opcode_type, 16#10#),
      2473 => to_slv(opcode_type, 16#09#),
      2474 => to_slv(opcode_type, 16#11#),
      2475 => to_slv(opcode_type, 16#0B#),
      2476 => to_slv(opcode_type, 16#06#),
      2477 => to_slv(opcode_type, 16#08#),
      2478 => to_slv(opcode_type, 16#0B#),
      2479 => to_slv(opcode_type, 16#0F#),
      2480 => to_slv(opcode_type, 16#09#),
      2481 => to_slv(opcode_type, 16#0F#),
      2482 => to_slv(opcode_type, 16#0F#),
      2483 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#07#),
      2497 => to_slv(opcode_type, 16#09#),
      2498 => to_slv(opcode_type, 16#09#),
      2499 => to_slv(opcode_type, 16#01#),
      2500 => to_slv(opcode_type, 16#0F#),
      2501 => to_slv(opcode_type, 16#06#),
      2502 => to_slv(opcode_type, 16#0A#),
      2503 => to_slv(opcode_type, 16#0A#),
      2504 => to_slv(opcode_type, 16#08#),
      2505 => to_slv(opcode_type, 16#01#),
      2506 => to_slv(opcode_type, 16#0D#),
      2507 => to_slv(opcode_type, 16#02#),
      2508 => to_slv(opcode_type, 16#0D#),
      2509 => to_slv(opcode_type, 16#01#),
      2510 => to_slv(opcode_type, 16#06#),
      2511 => to_slv(opcode_type, 16#08#),
      2512 => to_slv(opcode_type, 16#0E#),
      2513 => to_slv(opcode_type, 16#0C#),
      2514 => to_slv(opcode_type, 16#10#),
      2515 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#05#),
      2530 => to_slv(opcode_type, 16#02#),
      2531 => to_slv(opcode_type, 16#08#),
      2532 => to_slv(opcode_type, 16#0D#),
      2533 => to_slv(opcode_type, 16#11#),
      2534 => to_slv(opcode_type, 16#09#),
      2535 => to_slv(opcode_type, 16#09#),
      2536 => to_slv(opcode_type, 16#09#),
      2537 => to_slv(opcode_type, 16#0F#),
      2538 => to_slv(opcode_type, 16#0B#),
      2539 => to_slv(opcode_type, 16#04#),
      2540 => to_slv(opcode_type, 16#0D#),
      2541 => to_slv(opcode_type, 16#09#),
      2542 => to_slv(opcode_type, 16#03#),
      2543 => to_slv(opcode_type, 16#0B#),
      2544 => to_slv(opcode_type, 16#06#),
      2545 => to_slv(opcode_type, 16#0F#),
      2546 => to_slv(opcode_type, 16#10#),
      2547 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#09#),
      2561 => to_slv(opcode_type, 16#06#),
      2562 => to_slv(opcode_type, 16#08#),
      2563 => to_slv(opcode_type, 16#06#),
      2564 => to_slv(opcode_type, 16#0A#),
      2565 => to_slv(opcode_type, 16#11#),
      2566 => to_slv(opcode_type, 16#04#),
      2567 => to_slv(opcode_type, 16#10#),
      2568 => to_slv(opcode_type, 16#07#),
      2569 => to_slv(opcode_type, 16#07#),
      2570 => to_slv(opcode_type, 16#0B#),
      2571 => to_slv(opcode_type, 16#0D#),
      2572 => to_slv(opcode_type, 16#08#),
      2573 => to_slv(opcode_type, 16#0E#),
      2574 => to_slv(opcode_type, 16#0B#),
      2575 => to_slv(opcode_type, 16#07#),
      2576 => to_slv(opcode_type, 16#04#),
      2577 => to_slv(opcode_type, 16#0D#),
      2578 => to_slv(opcode_type, 16#0B#),
      2579 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#09#),
      2593 => to_slv(opcode_type, 16#08#),
      2594 => to_slv(opcode_type, 16#05#),
      2595 => to_slv(opcode_type, 16#01#),
      2596 => to_slv(opcode_type, 16#11#),
      2597 => to_slv(opcode_type, 16#02#),
      2598 => to_slv(opcode_type, 16#08#),
      2599 => to_slv(opcode_type, 16#B2#),
      2600 => to_slv(opcode_type, 16#0E#),
      2601 => to_slv(opcode_type, 16#07#),
      2602 => to_slv(opcode_type, 16#02#),
      2603 => to_slv(opcode_type, 16#02#),
      2604 => to_slv(opcode_type, 16#0D#),
      2605 => to_slv(opcode_type, 16#06#),
      2606 => to_slv(opcode_type, 16#08#),
      2607 => to_slv(opcode_type, 16#E8#),
      2608 => to_slv(opcode_type, 16#10#),
      2609 => to_slv(opcode_type, 16#03#),
      2610 => to_slv(opcode_type, 16#47#),
      2611 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#06#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#01#),
      2627 => to_slv(opcode_type, 16#01#),
      2628 => to_slv(opcode_type, 16#10#),
      2629 => to_slv(opcode_type, 16#06#),
      2630 => to_slv(opcode_type, 16#02#),
      2631 => to_slv(opcode_type, 16#0D#),
      2632 => to_slv(opcode_type, 16#04#),
      2633 => to_slv(opcode_type, 16#0C#),
      2634 => to_slv(opcode_type, 16#07#),
      2635 => to_slv(opcode_type, 16#09#),
      2636 => to_slv(opcode_type, 16#03#),
      2637 => to_slv(opcode_type, 16#0C#),
      2638 => to_slv(opcode_type, 16#03#),
      2639 => to_slv(opcode_type, 16#0C#),
      2640 => to_slv(opcode_type, 16#07#),
      2641 => to_slv(opcode_type, 16#0D#),
      2642 => to_slv(opcode_type, 16#0A#),
      2643 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#06#),
      2657 => to_slv(opcode_type, 16#09#),
      2658 => to_slv(opcode_type, 16#04#),
      2659 => to_slv(opcode_type, 16#08#),
      2660 => to_slv(opcode_type, 16#0E#),
      2661 => to_slv(opcode_type, 16#0F#),
      2662 => to_slv(opcode_type, 16#01#),
      2663 => to_slv(opcode_type, 16#02#),
      2664 => to_slv(opcode_type, 16#0E#),
      2665 => to_slv(opcode_type, 16#08#),
      2666 => to_slv(opcode_type, 16#01#),
      2667 => to_slv(opcode_type, 16#09#),
      2668 => to_slv(opcode_type, 16#10#),
      2669 => to_slv(opcode_type, 16#0A#),
      2670 => to_slv(opcode_type, 16#08#),
      2671 => to_slv(opcode_type, 16#09#),
      2672 => to_slv(opcode_type, 16#0D#),
      2673 => to_slv(opcode_type, 16#0A#),
      2674 => to_slv(opcode_type, 16#0E#),
      2675 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#09#),
      2689 => to_slv(opcode_type, 16#07#),
      2690 => to_slv(opcode_type, 16#07#),
      2691 => to_slv(opcode_type, 16#08#),
      2692 => to_slv(opcode_type, 16#10#),
      2693 => to_slv(opcode_type, 16#11#),
      2694 => to_slv(opcode_type, 16#07#),
      2695 => to_slv(opcode_type, 16#0D#),
      2696 => to_slv(opcode_type, 16#0A#),
      2697 => to_slv(opcode_type, 16#08#),
      2698 => to_slv(opcode_type, 16#04#),
      2699 => to_slv(opcode_type, 16#0E#),
      2700 => to_slv(opcode_type, 16#01#),
      2701 => to_slv(opcode_type, 16#0A#),
      2702 => to_slv(opcode_type, 16#06#),
      2703 => to_slv(opcode_type, 16#01#),
      2704 => to_slv(opcode_type, 16#02#),
      2705 => to_slv(opcode_type, 16#0F#),
      2706 => to_slv(opcode_type, 16#10#),
      2707 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#07#),
      2721 => to_slv(opcode_type, 16#02#),
      2722 => to_slv(opcode_type, 16#08#),
      2723 => to_slv(opcode_type, 16#08#),
      2724 => to_slv(opcode_type, 16#11#),
      2725 => to_slv(opcode_type, 16#0F#),
      2726 => to_slv(opcode_type, 16#04#),
      2727 => to_slv(opcode_type, 16#0A#),
      2728 => to_slv(opcode_type, 16#08#),
      2729 => to_slv(opcode_type, 16#02#),
      2730 => to_slv(opcode_type, 16#05#),
      2731 => to_slv(opcode_type, 16#25#),
      2732 => to_slv(opcode_type, 16#07#),
      2733 => to_slv(opcode_type, 16#07#),
      2734 => to_slv(opcode_type, 16#10#),
      2735 => to_slv(opcode_type, 16#0B#),
      2736 => to_slv(opcode_type, 16#09#),
      2737 => to_slv(opcode_type, 16#11#),
      2738 => to_slv(opcode_type, 16#0F#),
      2739 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#06#),
      2753 => to_slv(opcode_type, 16#01#),
      2754 => to_slv(opcode_type, 16#03#),
      2755 => to_slv(opcode_type, 16#09#),
      2756 => to_slv(opcode_type, 16#0C#),
      2757 => to_slv(opcode_type, 16#0F#),
      2758 => to_slv(opcode_type, 16#09#),
      2759 => to_slv(opcode_type, 16#09#),
      2760 => to_slv(opcode_type, 16#01#),
      2761 => to_slv(opcode_type, 16#DF#),
      2762 => to_slv(opcode_type, 16#03#),
      2763 => to_slv(opcode_type, 16#5B#),
      2764 => to_slv(opcode_type, 16#09#),
      2765 => to_slv(opcode_type, 16#09#),
      2766 => to_slv(opcode_type, 16#8A#),
      2767 => to_slv(opcode_type, 16#0B#),
      2768 => to_slv(opcode_type, 16#07#),
      2769 => to_slv(opcode_type, 16#0F#),
      2770 => to_slv(opcode_type, 16#0E#),
      2771 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#07#),
      2785 => to_slv(opcode_type, 16#04#),
      2786 => to_slv(opcode_type, 16#07#),
      2787 => to_slv(opcode_type, 16#03#),
      2788 => to_slv(opcode_type, 16#10#),
      2789 => to_slv(opcode_type, 16#06#),
      2790 => to_slv(opcode_type, 16#0E#),
      2791 => to_slv(opcode_type, 16#0C#),
      2792 => to_slv(opcode_type, 16#06#),
      2793 => to_slv(opcode_type, 16#09#),
      2794 => to_slv(opcode_type, 16#07#),
      2795 => to_slv(opcode_type, 16#11#),
      2796 => to_slv(opcode_type, 16#0C#),
      2797 => to_slv(opcode_type, 16#03#),
      2798 => to_slv(opcode_type, 16#0E#),
      2799 => to_slv(opcode_type, 16#07#),
      2800 => to_slv(opcode_type, 16#04#),
      2801 => to_slv(opcode_type, 16#10#),
      2802 => to_slv(opcode_type, 16#0C#),
      2803 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#08#),
      2817 => to_slv(opcode_type, 16#04#),
      2818 => to_slv(opcode_type, 16#08#),
      2819 => to_slv(opcode_type, 16#04#),
      2820 => to_slv(opcode_type, 16#11#),
      2821 => to_slv(opcode_type, 16#02#),
      2822 => to_slv(opcode_type, 16#0E#),
      2823 => to_slv(opcode_type, 16#08#),
      2824 => to_slv(opcode_type, 16#04#),
      2825 => to_slv(opcode_type, 16#09#),
      2826 => to_slv(opcode_type, 16#11#),
      2827 => to_slv(opcode_type, 16#10#),
      2828 => to_slv(opcode_type, 16#08#),
      2829 => to_slv(opcode_type, 16#08#),
      2830 => to_slv(opcode_type, 16#0A#),
      2831 => to_slv(opcode_type, 16#0C#),
      2832 => to_slv(opcode_type, 16#06#),
      2833 => to_slv(opcode_type, 16#0F#),
      2834 => to_slv(opcode_type, 16#0F#),
      2835 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#06#),
      2849 => to_slv(opcode_type, 16#02#),
      2850 => to_slv(opcode_type, 16#07#),
      2851 => to_slv(opcode_type, 16#01#),
      2852 => to_slv(opcode_type, 16#0F#),
      2853 => to_slv(opcode_type, 16#02#),
      2854 => to_slv(opcode_type, 16#0A#),
      2855 => to_slv(opcode_type, 16#08#),
      2856 => to_slv(opcode_type, 16#05#),
      2857 => to_slv(opcode_type, 16#06#),
      2858 => to_slv(opcode_type, 16#10#),
      2859 => to_slv(opcode_type, 16#0F#),
      2860 => to_slv(opcode_type, 16#08#),
      2861 => to_slv(opcode_type, 16#09#),
      2862 => to_slv(opcode_type, 16#0E#),
      2863 => to_slv(opcode_type, 16#0F#),
      2864 => to_slv(opcode_type, 16#08#),
      2865 => to_slv(opcode_type, 16#10#),
      2866 => to_slv(opcode_type, 16#0F#),
      2867 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#08#),
      2881 => to_slv(opcode_type, 16#04#),
      2882 => to_slv(opcode_type, 16#03#),
      2883 => to_slv(opcode_type, 16#08#),
      2884 => to_slv(opcode_type, 16#0C#),
      2885 => to_slv(opcode_type, 16#0C#),
      2886 => to_slv(opcode_type, 16#07#),
      2887 => to_slv(opcode_type, 16#06#),
      2888 => to_slv(opcode_type, 16#07#),
      2889 => to_slv(opcode_type, 16#0A#),
      2890 => to_slv(opcode_type, 16#0D#),
      2891 => to_slv(opcode_type, 16#01#),
      2892 => to_slv(opcode_type, 16#0C#),
      2893 => to_slv(opcode_type, 16#09#),
      2894 => to_slv(opcode_type, 16#01#),
      2895 => to_slv(opcode_type, 16#0D#),
      2896 => to_slv(opcode_type, 16#06#),
      2897 => to_slv(opcode_type, 16#0C#),
      2898 => to_slv(opcode_type, 16#0D#),
      2899 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#06#),
      2913 => to_slv(opcode_type, 16#08#),
      2914 => to_slv(opcode_type, 16#05#),
      2915 => to_slv(opcode_type, 16#09#),
      2916 => to_slv(opcode_type, 16#0F#),
      2917 => to_slv(opcode_type, 16#57#),
      2918 => to_slv(opcode_type, 16#08#),
      2919 => to_slv(opcode_type, 16#01#),
      2920 => to_slv(opcode_type, 16#0A#),
      2921 => to_slv(opcode_type, 16#06#),
      2922 => to_slv(opcode_type, 16#10#),
      2923 => to_slv(opcode_type, 16#0D#),
      2924 => to_slv(opcode_type, 16#05#),
      2925 => to_slv(opcode_type, 16#06#),
      2926 => to_slv(opcode_type, 16#06#),
      2927 => to_slv(opcode_type, 16#10#),
      2928 => to_slv(opcode_type, 16#10#),
      2929 => to_slv(opcode_type, 16#01#),
      2930 => to_slv(opcode_type, 16#0F#),
      2931 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#09#),
      2945 => to_slv(opcode_type, 16#09#),
      2946 => to_slv(opcode_type, 16#09#),
      2947 => to_slv(opcode_type, 16#06#),
      2948 => to_slv(opcode_type, 16#0D#),
      2949 => to_slv(opcode_type, 16#11#),
      2950 => to_slv(opcode_type, 16#02#),
      2951 => to_slv(opcode_type, 16#0A#),
      2952 => to_slv(opcode_type, 16#02#),
      2953 => to_slv(opcode_type, 16#07#),
      2954 => to_slv(opcode_type, 16#0B#),
      2955 => to_slv(opcode_type, 16#0D#),
      2956 => to_slv(opcode_type, 16#04#),
      2957 => to_slv(opcode_type, 16#09#),
      2958 => to_slv(opcode_type, 16#04#),
      2959 => to_slv(opcode_type, 16#11#),
      2960 => to_slv(opcode_type, 16#06#),
      2961 => to_slv(opcode_type, 16#0E#),
      2962 => to_slv(opcode_type, 16#11#),
      2963 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#06#),
      2977 => to_slv(opcode_type, 16#01#),
      2978 => to_slv(opcode_type, 16#03#),
      2979 => to_slv(opcode_type, 16#03#),
      2980 => to_slv(opcode_type, 16#D3#),
      2981 => to_slv(opcode_type, 16#07#),
      2982 => to_slv(opcode_type, 16#07#),
      2983 => to_slv(opcode_type, 16#04#),
      2984 => to_slv(opcode_type, 16#0E#),
      2985 => to_slv(opcode_type, 16#09#),
      2986 => to_slv(opcode_type, 16#AD#),
      2987 => to_slv(opcode_type, 16#0D#),
      2988 => to_slv(opcode_type, 16#08#),
      2989 => to_slv(opcode_type, 16#06#),
      2990 => to_slv(opcode_type, 16#0B#),
      2991 => to_slv(opcode_type, 16#0A#),
      2992 => to_slv(opcode_type, 16#09#),
      2993 => to_slv(opcode_type, 16#11#),
      2994 => to_slv(opcode_type, 16#10#),
      2995 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#07#),
      3009 => to_slv(opcode_type, 16#06#),
      3010 => to_slv(opcode_type, 16#01#),
      3011 => to_slv(opcode_type, 16#03#),
      3012 => to_slv(opcode_type, 16#0F#),
      3013 => to_slv(opcode_type, 16#01#),
      3014 => to_slv(opcode_type, 16#06#),
      3015 => to_slv(opcode_type, 16#10#),
      3016 => to_slv(opcode_type, 16#0B#),
      3017 => to_slv(opcode_type, 16#07#),
      3018 => to_slv(opcode_type, 16#09#),
      3019 => to_slv(opcode_type, 16#01#),
      3020 => to_slv(opcode_type, 16#0D#),
      3021 => to_slv(opcode_type, 16#01#),
      3022 => to_slv(opcode_type, 16#11#),
      3023 => to_slv(opcode_type, 16#03#),
      3024 => to_slv(opcode_type, 16#08#),
      3025 => to_slv(opcode_type, 16#0D#),
      3026 => to_slv(opcode_type, 16#0C#),
      3027 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#07#),
      3041 => to_slv(opcode_type, 16#01#),
      3042 => to_slv(opcode_type, 16#01#),
      3043 => to_slv(opcode_type, 16#03#),
      3044 => to_slv(opcode_type, 16#10#),
      3045 => to_slv(opcode_type, 16#09#),
      3046 => to_slv(opcode_type, 16#08#),
      3047 => to_slv(opcode_type, 16#09#),
      3048 => to_slv(opcode_type, 16#0D#),
      3049 => to_slv(opcode_type, 16#0D#),
      3050 => to_slv(opcode_type, 16#04#),
      3051 => to_slv(opcode_type, 16#0B#),
      3052 => to_slv(opcode_type, 16#09#),
      3053 => to_slv(opcode_type, 16#07#),
      3054 => to_slv(opcode_type, 16#0E#),
      3055 => to_slv(opcode_type, 16#0A#),
      3056 => to_slv(opcode_type, 16#07#),
      3057 => to_slv(opcode_type, 16#0A#),
      3058 => to_slv(opcode_type, 16#65#),
      3059 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#09#),
      3073 => to_slv(opcode_type, 16#08#),
      3074 => to_slv(opcode_type, 16#02#),
      3075 => to_slv(opcode_type, 16#08#),
      3076 => to_slv(opcode_type, 16#11#),
      3077 => to_slv(opcode_type, 16#0B#),
      3078 => to_slv(opcode_type, 16#05#),
      3079 => to_slv(opcode_type, 16#01#),
      3080 => to_slv(opcode_type, 16#84#),
      3081 => to_slv(opcode_type, 16#06#),
      3082 => to_slv(opcode_type, 16#02#),
      3083 => to_slv(opcode_type, 16#02#),
      3084 => to_slv(opcode_type, 16#0C#),
      3085 => to_slv(opcode_type, 16#09#),
      3086 => to_slv(opcode_type, 16#08#),
      3087 => to_slv(opcode_type, 16#0C#),
      3088 => to_slv(opcode_type, 16#0F#),
      3089 => to_slv(opcode_type, 16#03#),
      3090 => to_slv(opcode_type, 16#0C#),
      3091 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#06#),
      3105 => to_slv(opcode_type, 16#02#),
      3106 => to_slv(opcode_type, 16#01#),
      3107 => to_slv(opcode_type, 16#03#),
      3108 => to_slv(opcode_type, 16#52#),
      3109 => to_slv(opcode_type, 16#06#),
      3110 => to_slv(opcode_type, 16#08#),
      3111 => to_slv(opcode_type, 16#03#),
      3112 => to_slv(opcode_type, 16#43#),
      3113 => to_slv(opcode_type, 16#08#),
      3114 => to_slv(opcode_type, 16#10#),
      3115 => to_slv(opcode_type, 16#0A#),
      3116 => to_slv(opcode_type, 16#07#),
      3117 => to_slv(opcode_type, 16#08#),
      3118 => to_slv(opcode_type, 16#11#),
      3119 => to_slv(opcode_type, 16#0B#),
      3120 => to_slv(opcode_type, 16#09#),
      3121 => to_slv(opcode_type, 16#0B#),
      3122 => to_slv(opcode_type, 16#10#),
      3123 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#08#),
      3137 => to_slv(opcode_type, 16#09#),
      3138 => to_slv(opcode_type, 16#02#),
      3139 => to_slv(opcode_type, 16#06#),
      3140 => to_slv(opcode_type, 16#11#),
      3141 => to_slv(opcode_type, 16#10#),
      3142 => to_slv(opcode_type, 16#03#),
      3143 => to_slv(opcode_type, 16#05#),
      3144 => to_slv(opcode_type, 16#0C#),
      3145 => to_slv(opcode_type, 16#06#),
      3146 => to_slv(opcode_type, 16#06#),
      3147 => to_slv(opcode_type, 16#02#),
      3148 => to_slv(opcode_type, 16#13#),
      3149 => to_slv(opcode_type, 16#07#),
      3150 => to_slv(opcode_type, 16#0E#),
      3151 => to_slv(opcode_type, 16#11#),
      3152 => to_slv(opcode_type, 16#07#),
      3153 => to_slv(opcode_type, 16#0F#),
      3154 => to_slv(opcode_type, 16#11#),
      3155 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#06#),
      3169 => to_slv(opcode_type, 16#08#),
      3170 => to_slv(opcode_type, 16#04#),
      3171 => to_slv(opcode_type, 16#08#),
      3172 => to_slv(opcode_type, 16#0C#),
      3173 => to_slv(opcode_type, 16#52#),
      3174 => to_slv(opcode_type, 16#03#),
      3175 => to_slv(opcode_type, 16#02#),
      3176 => to_slv(opcode_type, 16#0A#),
      3177 => to_slv(opcode_type, 16#09#),
      3178 => to_slv(opcode_type, 16#07#),
      3179 => to_slv(opcode_type, 16#08#),
      3180 => to_slv(opcode_type, 16#0E#),
      3181 => to_slv(opcode_type, 16#0D#),
      3182 => to_slv(opcode_type, 16#04#),
      3183 => to_slv(opcode_type, 16#0A#),
      3184 => to_slv(opcode_type, 16#01#),
      3185 => to_slv(opcode_type, 16#04#),
      3186 => to_slv(opcode_type, 16#0C#),
      3187 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#06#),
      3201 => to_slv(opcode_type, 16#03#),
      3202 => to_slv(opcode_type, 16#06#),
      3203 => to_slv(opcode_type, 16#07#),
      3204 => to_slv(opcode_type, 16#10#),
      3205 => to_slv(opcode_type, 16#0D#),
      3206 => to_slv(opcode_type, 16#01#),
      3207 => to_slv(opcode_type, 16#10#),
      3208 => to_slv(opcode_type, 16#09#),
      3209 => to_slv(opcode_type, 16#01#),
      3210 => to_slv(opcode_type, 16#02#),
      3211 => to_slv(opcode_type, 16#0F#),
      3212 => to_slv(opcode_type, 16#06#),
      3213 => to_slv(opcode_type, 16#08#),
      3214 => to_slv(opcode_type, 16#11#),
      3215 => to_slv(opcode_type, 16#11#),
      3216 => to_slv(opcode_type, 16#08#),
      3217 => to_slv(opcode_type, 16#0B#),
      3218 => to_slv(opcode_type, 16#0E#),
      3219 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#08#),
      3233 => to_slv(opcode_type, 16#02#),
      3234 => to_slv(opcode_type, 16#06#),
      3235 => to_slv(opcode_type, 16#09#),
      3236 => to_slv(opcode_type, 16#10#),
      3237 => to_slv(opcode_type, 16#10#),
      3238 => to_slv(opcode_type, 16#02#),
      3239 => to_slv(opcode_type, 16#0A#),
      3240 => to_slv(opcode_type, 16#08#),
      3241 => to_slv(opcode_type, 16#04#),
      3242 => to_slv(opcode_type, 16#02#),
      3243 => to_slv(opcode_type, 16#0B#),
      3244 => to_slv(opcode_type, 16#08#),
      3245 => to_slv(opcode_type, 16#09#),
      3246 => to_slv(opcode_type, 16#0F#),
      3247 => to_slv(opcode_type, 16#0B#),
      3248 => to_slv(opcode_type, 16#06#),
      3249 => to_slv(opcode_type, 16#0A#),
      3250 => to_slv(opcode_type, 16#0E#),
      3251 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#07#),
      3265 => to_slv(opcode_type, 16#03#),
      3266 => to_slv(opcode_type, 16#06#),
      3267 => to_slv(opcode_type, 16#03#),
      3268 => to_slv(opcode_type, 16#11#),
      3269 => to_slv(opcode_type, 16#01#),
      3270 => to_slv(opcode_type, 16#10#),
      3271 => to_slv(opcode_type, 16#06#),
      3272 => to_slv(opcode_type, 16#04#),
      3273 => to_slv(opcode_type, 16#08#),
      3274 => to_slv(opcode_type, 16#10#),
      3275 => to_slv(opcode_type, 16#0A#),
      3276 => to_slv(opcode_type, 16#09#),
      3277 => to_slv(opcode_type, 16#08#),
      3278 => to_slv(opcode_type, 16#0D#),
      3279 => to_slv(opcode_type, 16#7B#),
      3280 => to_slv(opcode_type, 16#09#),
      3281 => to_slv(opcode_type, 16#0A#),
      3282 => to_slv(opcode_type, 16#0C#),
      3283 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#09#),
      3297 => to_slv(opcode_type, 16#01#),
      3298 => to_slv(opcode_type, 16#04#),
      3299 => to_slv(opcode_type, 16#01#),
      3300 => to_slv(opcode_type, 16#AE#),
      3301 => to_slv(opcode_type, 16#09#),
      3302 => to_slv(opcode_type, 16#06#),
      3303 => to_slv(opcode_type, 16#08#),
      3304 => to_slv(opcode_type, 16#AF#),
      3305 => to_slv(opcode_type, 16#0E#),
      3306 => to_slv(opcode_type, 16#04#),
      3307 => to_slv(opcode_type, 16#10#),
      3308 => to_slv(opcode_type, 16#09#),
      3309 => to_slv(opcode_type, 16#07#),
      3310 => to_slv(opcode_type, 16#10#),
      3311 => to_slv(opcode_type, 16#11#),
      3312 => to_slv(opcode_type, 16#06#),
      3313 => to_slv(opcode_type, 16#0F#),
      3314 => to_slv(opcode_type, 16#56#),
      3315 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#09#),
      3329 => to_slv(opcode_type, 16#04#),
      3330 => to_slv(opcode_type, 16#05#),
      3331 => to_slv(opcode_type, 16#02#),
      3332 => to_slv(opcode_type, 16#45#),
      3333 => to_slv(opcode_type, 16#07#),
      3334 => to_slv(opcode_type, 16#08#),
      3335 => to_slv(opcode_type, 16#08#),
      3336 => to_slv(opcode_type, 16#B1#),
      3337 => to_slv(opcode_type, 16#23#),
      3338 => to_slv(opcode_type, 16#07#),
      3339 => to_slv(opcode_type, 16#68#),
      3340 => to_slv(opcode_type, 16#10#),
      3341 => to_slv(opcode_type, 16#07#),
      3342 => to_slv(opcode_type, 16#09#),
      3343 => to_slv(opcode_type, 16#3F#),
      3344 => to_slv(opcode_type, 16#0D#),
      3345 => to_slv(opcode_type, 16#05#),
      3346 => to_slv(opcode_type, 16#0D#),
      3347 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#07#),
      3361 => to_slv(opcode_type, 16#02#),
      3362 => to_slv(opcode_type, 16#03#),
      3363 => to_slv(opcode_type, 16#03#),
      3364 => to_slv(opcode_type, 16#E9#),
      3365 => to_slv(opcode_type, 16#06#),
      3366 => to_slv(opcode_type, 16#07#),
      3367 => to_slv(opcode_type, 16#01#),
      3368 => to_slv(opcode_type, 16#0F#),
      3369 => to_slv(opcode_type, 16#06#),
      3370 => to_slv(opcode_type, 16#0C#),
      3371 => to_slv(opcode_type, 16#0F#),
      3372 => to_slv(opcode_type, 16#06#),
      3373 => to_slv(opcode_type, 16#08#),
      3374 => to_slv(opcode_type, 16#0E#),
      3375 => to_slv(opcode_type, 16#0B#),
      3376 => to_slv(opcode_type, 16#09#),
      3377 => to_slv(opcode_type, 16#0B#),
      3378 => to_slv(opcode_type, 16#0D#),
      3379 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#08#),
      3393 => to_slv(opcode_type, 16#07#),
      3394 => to_slv(opcode_type, 16#01#),
      3395 => to_slv(opcode_type, 16#02#),
      3396 => to_slv(opcode_type, 16#93#),
      3397 => to_slv(opcode_type, 16#04#),
      3398 => to_slv(opcode_type, 16#06#),
      3399 => to_slv(opcode_type, 16#0C#),
      3400 => to_slv(opcode_type, 16#0B#),
      3401 => to_slv(opcode_type, 16#06#),
      3402 => to_slv(opcode_type, 16#03#),
      3403 => to_slv(opcode_type, 16#06#),
      3404 => to_slv(opcode_type, 16#0F#),
      3405 => to_slv(opcode_type, 16#0E#),
      3406 => to_slv(opcode_type, 16#08#),
      3407 => to_slv(opcode_type, 16#03#),
      3408 => to_slv(opcode_type, 16#0F#),
      3409 => to_slv(opcode_type, 16#05#),
      3410 => to_slv(opcode_type, 16#0A#),
      3411 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#08#),
      3426 => to_slv(opcode_type, 16#08#),
      3427 => to_slv(opcode_type, 16#05#),
      3428 => to_slv(opcode_type, 16#1F#),
      3429 => to_slv(opcode_type, 16#04#),
      3430 => to_slv(opcode_type, 16#0B#),
      3431 => to_slv(opcode_type, 16#01#),
      3432 => to_slv(opcode_type, 16#03#),
      3433 => to_slv(opcode_type, 16#0E#),
      3434 => to_slv(opcode_type, 16#09#),
      3435 => to_slv(opcode_type, 16#03#),
      3436 => to_slv(opcode_type, 16#09#),
      3437 => to_slv(opcode_type, 16#10#),
      3438 => to_slv(opcode_type, 16#11#),
      3439 => to_slv(opcode_type, 16#01#),
      3440 => to_slv(opcode_type, 16#09#),
      3441 => to_slv(opcode_type, 16#0A#),
      3442 => to_slv(opcode_type, 16#0E#),
      3443 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#06#),
      3457 => to_slv(opcode_type, 16#09#),
      3458 => to_slv(opcode_type, 16#07#),
      3459 => to_slv(opcode_type, 16#04#),
      3460 => to_slv(opcode_type, 16#11#),
      3461 => to_slv(opcode_type, 16#06#),
      3462 => to_slv(opcode_type, 16#0E#),
      3463 => to_slv(opcode_type, 16#85#),
      3464 => to_slv(opcode_type, 16#02#),
      3465 => to_slv(opcode_type, 16#06#),
      3466 => to_slv(opcode_type, 16#D5#),
      3467 => to_slv(opcode_type, 16#0D#),
      3468 => to_slv(opcode_type, 16#05#),
      3469 => to_slv(opcode_type, 16#09#),
      3470 => to_slv(opcode_type, 16#07#),
      3471 => to_slv(opcode_type, 16#0B#),
      3472 => to_slv(opcode_type, 16#46#),
      3473 => to_slv(opcode_type, 16#02#),
      3474 => to_slv(opcode_type, 16#10#),
      3475 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#07#),
      3489 => to_slv(opcode_type, 16#01#),
      3490 => to_slv(opcode_type, 16#08#),
      3491 => to_slv(opcode_type, 16#08#),
      3492 => to_slv(opcode_type, 16#0A#),
      3493 => to_slv(opcode_type, 16#0D#),
      3494 => to_slv(opcode_type, 16#06#),
      3495 => to_slv(opcode_type, 16#0E#),
      3496 => to_slv(opcode_type, 16#F0#),
      3497 => to_slv(opcode_type, 16#06#),
      3498 => to_slv(opcode_type, 16#04#),
      3499 => to_slv(opcode_type, 16#06#),
      3500 => to_slv(opcode_type, 16#0A#),
      3501 => to_slv(opcode_type, 16#0C#),
      3502 => to_slv(opcode_type, 16#08#),
      3503 => to_slv(opcode_type, 16#04#),
      3504 => to_slv(opcode_type, 16#10#),
      3505 => to_slv(opcode_type, 16#04#),
      3506 => to_slv(opcode_type, 16#0D#),
      3507 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#09#),
      3521 => to_slv(opcode_type, 16#03#),
      3522 => to_slv(opcode_type, 16#03#),
      3523 => to_slv(opcode_type, 16#09#),
      3524 => to_slv(opcode_type, 16#10#),
      3525 => to_slv(opcode_type, 16#0F#),
      3526 => to_slv(opcode_type, 16#06#),
      3527 => to_slv(opcode_type, 16#08#),
      3528 => to_slv(opcode_type, 16#03#),
      3529 => to_slv(opcode_type, 16#11#),
      3530 => to_slv(opcode_type, 16#07#),
      3531 => to_slv(opcode_type, 16#10#),
      3532 => to_slv(opcode_type, 16#0B#),
      3533 => to_slv(opcode_type, 16#06#),
      3534 => to_slv(opcode_type, 16#04#),
      3535 => to_slv(opcode_type, 16#0E#),
      3536 => to_slv(opcode_type, 16#08#),
      3537 => to_slv(opcode_type, 16#0D#),
      3538 => to_slv(opcode_type, 16#0B#),
      3539 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#07#),
      3553 => to_slv(opcode_type, 16#08#),
      3554 => to_slv(opcode_type, 16#08#),
      3555 => to_slv(opcode_type, 16#04#),
      3556 => to_slv(opcode_type, 16#10#),
      3557 => to_slv(opcode_type, 16#07#),
      3558 => to_slv(opcode_type, 16#0B#),
      3559 => to_slv(opcode_type, 16#0C#),
      3560 => to_slv(opcode_type, 16#07#),
      3561 => to_slv(opcode_type, 16#01#),
      3562 => to_slv(opcode_type, 16#0D#),
      3563 => to_slv(opcode_type, 16#02#),
      3564 => to_slv(opcode_type, 16#0C#),
      3565 => to_slv(opcode_type, 16#04#),
      3566 => to_slv(opcode_type, 16#07#),
      3567 => to_slv(opcode_type, 16#09#),
      3568 => to_slv(opcode_type, 16#0E#),
      3569 => to_slv(opcode_type, 16#93#),
      3570 => to_slv(opcode_type, 16#0E#),
      3571 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#09#),
      3585 => to_slv(opcode_type, 16#08#),
      3586 => to_slv(opcode_type, 16#09#),
      3587 => to_slv(opcode_type, 16#08#),
      3588 => to_slv(opcode_type, 16#10#),
      3589 => to_slv(opcode_type, 16#10#),
      3590 => to_slv(opcode_type, 16#08#),
      3591 => to_slv(opcode_type, 16#10#),
      3592 => to_slv(opcode_type, 16#0B#),
      3593 => to_slv(opcode_type, 16#05#),
      3594 => to_slv(opcode_type, 16#07#),
      3595 => to_slv(opcode_type, 16#0B#),
      3596 => to_slv(opcode_type, 16#0A#),
      3597 => to_slv(opcode_type, 16#01#),
      3598 => to_slv(opcode_type, 16#06#),
      3599 => to_slv(opcode_type, 16#04#),
      3600 => to_slv(opcode_type, 16#0D#),
      3601 => to_slv(opcode_type, 16#01#),
      3602 => to_slv(opcode_type, 16#11#),
      3603 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#07#),
      3617 => to_slv(opcode_type, 16#06#),
      3618 => to_slv(opcode_type, 16#03#),
      3619 => to_slv(opcode_type, 16#09#),
      3620 => to_slv(opcode_type, 16#0E#),
      3621 => to_slv(opcode_type, 16#10#),
      3622 => to_slv(opcode_type, 16#05#),
      3623 => to_slv(opcode_type, 16#03#),
      3624 => to_slv(opcode_type, 16#0A#),
      3625 => to_slv(opcode_type, 16#09#),
      3626 => to_slv(opcode_type, 16#02#),
      3627 => to_slv(opcode_type, 16#05#),
      3628 => to_slv(opcode_type, 16#11#),
      3629 => to_slv(opcode_type, 16#08#),
      3630 => to_slv(opcode_type, 16#04#),
      3631 => to_slv(opcode_type, 16#10#),
      3632 => to_slv(opcode_type, 16#08#),
      3633 => to_slv(opcode_type, 16#0F#),
      3634 => to_slv(opcode_type, 16#0B#),
      3635 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#09#),
      3649 => to_slv(opcode_type, 16#08#),
      3650 => to_slv(opcode_type, 16#09#),
      3651 => to_slv(opcode_type, 16#01#),
      3652 => to_slv(opcode_type, 16#0A#),
      3653 => to_slv(opcode_type, 16#05#),
      3654 => to_slv(opcode_type, 16#0E#),
      3655 => to_slv(opcode_type, 16#06#),
      3656 => to_slv(opcode_type, 16#08#),
      3657 => to_slv(opcode_type, 16#0B#),
      3658 => to_slv(opcode_type, 16#11#),
      3659 => to_slv(opcode_type, 16#03#),
      3660 => to_slv(opcode_type, 16#0C#),
      3661 => to_slv(opcode_type, 16#08#),
      3662 => to_slv(opcode_type, 16#05#),
      3663 => to_slv(opcode_type, 16#04#),
      3664 => to_slv(opcode_type, 16#0F#),
      3665 => to_slv(opcode_type, 16#01#),
      3666 => to_slv(opcode_type, 16#0C#),
      3667 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#09#),
      3681 => to_slv(opcode_type, 16#07#),
      3682 => to_slv(opcode_type, 16#07#),
      3683 => to_slv(opcode_type, 16#04#),
      3684 => to_slv(opcode_type, 16#0C#),
      3685 => to_slv(opcode_type, 16#04#),
      3686 => to_slv(opcode_type, 16#0F#),
      3687 => to_slv(opcode_type, 16#02#),
      3688 => to_slv(opcode_type, 16#01#),
      3689 => to_slv(opcode_type, 16#0C#),
      3690 => to_slv(opcode_type, 16#08#),
      3691 => to_slv(opcode_type, 16#04#),
      3692 => to_slv(opcode_type, 16#02#),
      3693 => to_slv(opcode_type, 16#0A#),
      3694 => to_slv(opcode_type, 16#07#),
      3695 => to_slv(opcode_type, 16#05#),
      3696 => to_slv(opcode_type, 16#0A#),
      3697 => to_slv(opcode_type, 16#03#),
      3698 => to_slv(opcode_type, 16#0E#),
      3699 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#06#),
      3713 => to_slv(opcode_type, 16#01#),
      3714 => to_slv(opcode_type, 16#05#),
      3715 => to_slv(opcode_type, 16#07#),
      3716 => to_slv(opcode_type, 16#0A#),
      3717 => to_slv(opcode_type, 16#0B#),
      3718 => to_slv(opcode_type, 16#07#),
      3719 => to_slv(opcode_type, 16#08#),
      3720 => to_slv(opcode_type, 16#09#),
      3721 => to_slv(opcode_type, 16#CD#),
      3722 => to_slv(opcode_type, 16#10#),
      3723 => to_slv(opcode_type, 16#01#),
      3724 => to_slv(opcode_type, 16#0E#),
      3725 => to_slv(opcode_type, 16#09#),
      3726 => to_slv(opcode_type, 16#06#),
      3727 => to_slv(opcode_type, 16#0F#),
      3728 => to_slv(opcode_type, 16#0D#),
      3729 => to_slv(opcode_type, 16#03#),
      3730 => to_slv(opcode_type, 16#0C#),
      3731 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#08#),
      3745 => to_slv(opcode_type, 16#03#),
      3746 => to_slv(opcode_type, 16#02#),
      3747 => to_slv(opcode_type, 16#08#),
      3748 => to_slv(opcode_type, 16#FE#),
      3749 => to_slv(opcode_type, 16#0F#),
      3750 => to_slv(opcode_type, 16#08#),
      3751 => to_slv(opcode_type, 16#08#),
      3752 => to_slv(opcode_type, 16#06#),
      3753 => to_slv(opcode_type, 16#9F#),
      3754 => to_slv(opcode_type, 16#10#),
      3755 => to_slv(opcode_type, 16#05#),
      3756 => to_slv(opcode_type, 16#0D#),
      3757 => to_slv(opcode_type, 16#06#),
      3758 => to_slv(opcode_type, 16#07#),
      3759 => to_slv(opcode_type, 16#0F#),
      3760 => to_slv(opcode_type, 16#0B#),
      3761 => to_slv(opcode_type, 16#04#),
      3762 => to_slv(opcode_type, 16#0E#),
      3763 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#09#),
      3777 => to_slv(opcode_type, 16#07#),
      3778 => to_slv(opcode_type, 16#01#),
      3779 => to_slv(opcode_type, 16#05#),
      3780 => to_slv(opcode_type, 16#0D#),
      3781 => to_slv(opcode_type, 16#02#),
      3782 => to_slv(opcode_type, 16#03#),
      3783 => to_slv(opcode_type, 16#0B#),
      3784 => to_slv(opcode_type, 16#08#),
      3785 => to_slv(opcode_type, 16#02#),
      3786 => to_slv(opcode_type, 16#06#),
      3787 => to_slv(opcode_type, 16#0F#),
      3788 => to_slv(opcode_type, 16#24#),
      3789 => to_slv(opcode_type, 16#08#),
      3790 => to_slv(opcode_type, 16#01#),
      3791 => to_slv(opcode_type, 16#11#),
      3792 => to_slv(opcode_type, 16#08#),
      3793 => to_slv(opcode_type, 16#0F#),
      3794 => to_slv(opcode_type, 16#0E#),
      3795 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#08#),
      3809 => to_slv(opcode_type, 16#05#),
      3810 => to_slv(opcode_type, 16#05#),
      3811 => to_slv(opcode_type, 16#08#),
      3812 => to_slv(opcode_type, 16#0A#),
      3813 => to_slv(opcode_type, 16#0D#),
      3814 => to_slv(opcode_type, 16#08#),
      3815 => to_slv(opcode_type, 16#09#),
      3816 => to_slv(opcode_type, 16#02#),
      3817 => to_slv(opcode_type, 16#11#),
      3818 => to_slv(opcode_type, 16#04#),
      3819 => to_slv(opcode_type, 16#0D#),
      3820 => to_slv(opcode_type, 16#09#),
      3821 => to_slv(opcode_type, 16#09#),
      3822 => to_slv(opcode_type, 16#0B#),
      3823 => to_slv(opcode_type, 16#0B#),
      3824 => to_slv(opcode_type, 16#09#),
      3825 => to_slv(opcode_type, 16#0D#),
      3826 => to_slv(opcode_type, 16#10#),
      3827 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#08#),
      3841 => to_slv(opcode_type, 16#04#),
      3842 => to_slv(opcode_type, 16#09#),
      3843 => to_slv(opcode_type, 16#03#),
      3844 => to_slv(opcode_type, 16#B1#),
      3845 => to_slv(opcode_type, 16#04#),
      3846 => to_slv(opcode_type, 16#11#),
      3847 => to_slv(opcode_type, 16#09#),
      3848 => to_slv(opcode_type, 16#01#),
      3849 => to_slv(opcode_type, 16#06#),
      3850 => to_slv(opcode_type, 16#0A#),
      3851 => to_slv(opcode_type, 16#10#),
      3852 => to_slv(opcode_type, 16#08#),
      3853 => to_slv(opcode_type, 16#09#),
      3854 => to_slv(opcode_type, 16#0C#),
      3855 => to_slv(opcode_type, 16#0E#),
      3856 => to_slv(opcode_type, 16#09#),
      3857 => to_slv(opcode_type, 16#0F#),
      3858 => to_slv(opcode_type, 16#0F#),
      3859 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#09#),
      3873 => to_slv(opcode_type, 16#08#),
      3874 => to_slv(opcode_type, 16#03#),
      3875 => to_slv(opcode_type, 16#03#),
      3876 => to_slv(opcode_type, 16#0A#),
      3877 => to_slv(opcode_type, 16#08#),
      3878 => to_slv(opcode_type, 16#09#),
      3879 => to_slv(opcode_type, 16#0E#),
      3880 => to_slv(opcode_type, 16#70#),
      3881 => to_slv(opcode_type, 16#03#),
      3882 => to_slv(opcode_type, 16#E6#),
      3883 => to_slv(opcode_type, 16#03#),
      3884 => to_slv(opcode_type, 16#07#),
      3885 => to_slv(opcode_type, 16#09#),
      3886 => to_slv(opcode_type, 16#0E#),
      3887 => to_slv(opcode_type, 16#0E#),
      3888 => to_slv(opcode_type, 16#07#),
      3889 => to_slv(opcode_type, 16#0E#),
      3890 => to_slv(opcode_type, 16#11#),
      3891 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#08#),
      3905 => to_slv(opcode_type, 16#05#),
      3906 => to_slv(opcode_type, 16#02#),
      3907 => to_slv(opcode_type, 16#03#),
      3908 => to_slv(opcode_type, 16#10#),
      3909 => to_slv(opcode_type, 16#08#),
      3910 => to_slv(opcode_type, 16#08#),
      3911 => to_slv(opcode_type, 16#03#),
      3912 => to_slv(opcode_type, 16#41#),
      3913 => to_slv(opcode_type, 16#09#),
      3914 => to_slv(opcode_type, 16#11#),
      3915 => to_slv(opcode_type, 16#0E#),
      3916 => to_slv(opcode_type, 16#06#),
      3917 => to_slv(opcode_type, 16#06#),
      3918 => to_slv(opcode_type, 16#0A#),
      3919 => to_slv(opcode_type, 16#0D#),
      3920 => to_slv(opcode_type, 16#08#),
      3921 => to_slv(opcode_type, 16#11#),
      3922 => to_slv(opcode_type, 16#0F#),
      3923 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#06#),
      3937 => to_slv(opcode_type, 16#02#),
      3938 => to_slv(opcode_type, 16#02#),
      3939 => to_slv(opcode_type, 16#06#),
      3940 => to_slv(opcode_type, 16#0E#),
      3941 => to_slv(opcode_type, 16#10#),
      3942 => to_slv(opcode_type, 16#06#),
      3943 => to_slv(opcode_type, 16#08#),
      3944 => to_slv(opcode_type, 16#05#),
      3945 => to_slv(opcode_type, 16#0B#),
      3946 => to_slv(opcode_type, 16#01#),
      3947 => to_slv(opcode_type, 16#0B#),
      3948 => to_slv(opcode_type, 16#09#),
      3949 => to_slv(opcode_type, 16#08#),
      3950 => to_slv(opcode_type, 16#0A#),
      3951 => to_slv(opcode_type, 16#0C#),
      3952 => to_slv(opcode_type, 16#08#),
      3953 => to_slv(opcode_type, 16#0C#),
      3954 => to_slv(opcode_type, 16#0D#),
      3955 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#08#),
      3969 => to_slv(opcode_type, 16#01#),
      3970 => to_slv(opcode_type, 16#04#),
      3971 => to_slv(opcode_type, 16#03#),
      3972 => to_slv(opcode_type, 16#0B#),
      3973 => to_slv(opcode_type, 16#09#),
      3974 => to_slv(opcode_type, 16#06#),
      3975 => to_slv(opcode_type, 16#06#),
      3976 => to_slv(opcode_type, 16#0A#),
      3977 => to_slv(opcode_type, 16#0C#),
      3978 => to_slv(opcode_type, 16#05#),
      3979 => to_slv(opcode_type, 16#39#),
      3980 => to_slv(opcode_type, 16#09#),
      3981 => to_slv(opcode_type, 16#06#),
      3982 => to_slv(opcode_type, 16#0F#),
      3983 => to_slv(opcode_type, 16#0D#),
      3984 => to_slv(opcode_type, 16#08#),
      3985 => to_slv(opcode_type, 16#6E#),
      3986 => to_slv(opcode_type, 16#0E#),
      3987 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#08#),
      4001 => to_slv(opcode_type, 16#02#),
      4002 => to_slv(opcode_type, 16#04#),
      4003 => to_slv(opcode_type, 16#05#),
      4004 => to_slv(opcode_type, 16#10#),
      4005 => to_slv(opcode_type, 16#06#),
      4006 => to_slv(opcode_type, 16#08#),
      4007 => to_slv(opcode_type, 16#07#),
      4008 => to_slv(opcode_type, 16#11#),
      4009 => to_slv(opcode_type, 16#EA#),
      4010 => to_slv(opcode_type, 16#01#),
      4011 => to_slv(opcode_type, 16#11#),
      4012 => to_slv(opcode_type, 16#08#),
      4013 => to_slv(opcode_type, 16#06#),
      4014 => to_slv(opcode_type, 16#0F#),
      4015 => to_slv(opcode_type, 16#0F#),
      4016 => to_slv(opcode_type, 16#08#),
      4017 => to_slv(opcode_type, 16#10#),
      4018 => to_slv(opcode_type, 16#0E#),
      4019 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#07#),
      4033 => to_slv(opcode_type, 16#01#),
      4034 => to_slv(opcode_type, 16#04#),
      4035 => to_slv(opcode_type, 16#03#),
      4036 => to_slv(opcode_type, 16#0E#),
      4037 => to_slv(opcode_type, 16#06#),
      4038 => to_slv(opcode_type, 16#09#),
      4039 => to_slv(opcode_type, 16#04#),
      4040 => to_slv(opcode_type, 16#11#),
      4041 => to_slv(opcode_type, 16#09#),
      4042 => to_slv(opcode_type, 16#4D#),
      4043 => to_slv(opcode_type, 16#0D#),
      4044 => to_slv(opcode_type, 16#09#),
      4045 => to_slv(opcode_type, 16#08#),
      4046 => to_slv(opcode_type, 16#10#),
      4047 => to_slv(opcode_type, 16#0B#),
      4048 => to_slv(opcode_type, 16#08#),
      4049 => to_slv(opcode_type, 16#11#),
      4050 => to_slv(opcode_type, 16#0D#),
      4051 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#07#),
      4065 => to_slv(opcode_type, 16#09#),
      4066 => to_slv(opcode_type, 16#05#),
      4067 => to_slv(opcode_type, 16#09#),
      4068 => to_slv(opcode_type, 16#0D#),
      4069 => to_slv(opcode_type, 16#11#),
      4070 => to_slv(opcode_type, 16#04#),
      4071 => to_slv(opcode_type, 16#02#),
      4072 => to_slv(opcode_type, 16#3C#),
      4073 => to_slv(opcode_type, 16#06#),
      4074 => to_slv(opcode_type, 16#07#),
      4075 => to_slv(opcode_type, 16#03#),
      4076 => to_slv(opcode_type, 16#0A#),
      4077 => to_slv(opcode_type, 16#07#),
      4078 => to_slv(opcode_type, 16#0D#),
      4079 => to_slv(opcode_type, 16#0E#),
      4080 => to_slv(opcode_type, 16#04#),
      4081 => to_slv(opcode_type, 16#03#),
      4082 => to_slv(opcode_type, 16#10#),
      4083 to 4095 => (others => '0')
  ),

    -- Bin `20`...
    19 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#08#),
      1 => to_slv(opcode_type, 16#05#),
      2 => to_slv(opcode_type, 16#07#),
      3 => to_slv(opcode_type, 16#07#),
      4 => to_slv(opcode_type, 16#0C#),
      5 => to_slv(opcode_type, 16#0A#),
      6 => to_slv(opcode_type, 16#03#),
      7 => to_slv(opcode_type, 16#0F#),
      8 => to_slv(opcode_type, 16#08#),
      9 => to_slv(opcode_type, 16#06#),
      10 => to_slv(opcode_type, 16#08#),
      11 => to_slv(opcode_type, 16#0E#),
      12 => to_slv(opcode_type, 16#0C#),
      13 => to_slv(opcode_type, 16#05#),
      14 => to_slv(opcode_type, 16#0F#),
      15 => to_slv(opcode_type, 16#07#),
      16 => to_slv(opcode_type, 16#03#),
      17 => to_slv(opcode_type, 16#0B#),
      18 => to_slv(opcode_type, 16#05#),
      19 => to_slv(opcode_type, 16#9B#),
      20 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#09#),
      33 => to_slv(opcode_type, 16#07#),
      34 => to_slv(opcode_type, 16#06#),
      35 => to_slv(opcode_type, 16#09#),
      36 => to_slv(opcode_type, 16#0D#),
      37 => to_slv(opcode_type, 16#0E#),
      38 => to_slv(opcode_type, 16#04#),
      39 => to_slv(opcode_type, 16#11#),
      40 => to_slv(opcode_type, 16#05#),
      41 => to_slv(opcode_type, 16#04#),
      42 => to_slv(opcode_type, 16#0E#),
      43 => to_slv(opcode_type, 16#06#),
      44 => to_slv(opcode_type, 16#04#),
      45 => to_slv(opcode_type, 16#06#),
      46 => to_slv(opcode_type, 16#0D#),
      47 => to_slv(opcode_type, 16#0F#),
      48 => to_slv(opcode_type, 16#02#),
      49 => to_slv(opcode_type, 16#06#),
      50 => to_slv(opcode_type, 16#44#),
      51 => to_slv(opcode_type, 16#0C#),
      52 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#09#),
      65 => to_slv(opcode_type, 16#01#),
      66 => to_slv(opcode_type, 16#05#),
      67 => to_slv(opcode_type, 16#09#),
      68 => to_slv(opcode_type, 16#95#),
      69 => to_slv(opcode_type, 16#10#),
      70 => to_slv(opcode_type, 16#08#),
      71 => to_slv(opcode_type, 16#08#),
      72 => to_slv(opcode_type, 16#04#),
      73 => to_slv(opcode_type, 16#10#),
      74 => to_slv(opcode_type, 16#09#),
      75 => to_slv(opcode_type, 16#11#),
      76 => to_slv(opcode_type, 16#11#),
      77 => to_slv(opcode_type, 16#08#),
      78 => to_slv(opcode_type, 16#09#),
      79 => to_slv(opcode_type, 16#0B#),
      80 => to_slv(opcode_type, 16#0A#),
      81 => to_slv(opcode_type, 16#09#),
      82 => to_slv(opcode_type, 16#10#),
      83 => to_slv(opcode_type, 16#0E#),
      84 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#08#),
      97 => to_slv(opcode_type, 16#01#),
      98 => to_slv(opcode_type, 16#01#),
      99 => to_slv(opcode_type, 16#03#),
      100 => to_slv(opcode_type, 16#0A#),
      101 => to_slv(opcode_type, 16#09#),
      102 => to_slv(opcode_type, 16#09#),
      103 => to_slv(opcode_type, 16#09#),
      104 => to_slv(opcode_type, 16#0D#),
      105 => to_slv(opcode_type, 16#0A#),
      106 => to_slv(opcode_type, 16#07#),
      107 => to_slv(opcode_type, 16#0B#),
      108 => to_slv(opcode_type, 16#0C#),
      109 => to_slv(opcode_type, 16#09#),
      110 => to_slv(opcode_type, 16#08#),
      111 => to_slv(opcode_type, 16#0C#),
      112 => to_slv(opcode_type, 16#0D#),
      113 => to_slv(opcode_type, 16#06#),
      114 => to_slv(opcode_type, 16#0F#),
      115 => to_slv(opcode_type, 16#0D#),
      116 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#09#),
      129 => to_slv(opcode_type, 16#05#),
      130 => to_slv(opcode_type, 16#06#),
      131 => to_slv(opcode_type, 16#08#),
      132 => to_slv(opcode_type, 16#10#),
      133 => to_slv(opcode_type, 16#0D#),
      134 => to_slv(opcode_type, 16#04#),
      135 => to_slv(opcode_type, 16#0A#),
      136 => to_slv(opcode_type, 16#06#),
      137 => to_slv(opcode_type, 16#08#),
      138 => to_slv(opcode_type, 16#08#),
      139 => to_slv(opcode_type, 16#0D#),
      140 => to_slv(opcode_type, 16#0D#),
      141 => to_slv(opcode_type, 16#08#),
      142 => to_slv(opcode_type, 16#0A#),
      143 => to_slv(opcode_type, 16#0B#),
      144 => to_slv(opcode_type, 16#04#),
      145 => to_slv(opcode_type, 16#08#),
      146 => to_slv(opcode_type, 16#0F#),
      147 => to_slv(opcode_type, 16#0F#),
      148 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#07#),
      161 => to_slv(opcode_type, 16#04#),
      162 => to_slv(opcode_type, 16#04#),
      163 => to_slv(opcode_type, 16#01#),
      164 => to_slv(opcode_type, 16#D6#),
      165 => to_slv(opcode_type, 16#07#),
      166 => to_slv(opcode_type, 16#09#),
      167 => to_slv(opcode_type, 16#06#),
      168 => to_slv(opcode_type, 16#10#),
      169 => to_slv(opcode_type, 16#0A#),
      170 => to_slv(opcode_type, 16#06#),
      171 => to_slv(opcode_type, 16#10#),
      172 => to_slv(opcode_type, 16#0F#),
      173 => to_slv(opcode_type, 16#06#),
      174 => to_slv(opcode_type, 16#07#),
      175 => to_slv(opcode_type, 16#10#),
      176 => to_slv(opcode_type, 16#0D#),
      177 => to_slv(opcode_type, 16#06#),
      178 => to_slv(opcode_type, 16#0A#),
      179 => to_slv(opcode_type, 16#10#),
      180 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#08#),
      193 => to_slv(opcode_type, 16#02#),
      194 => to_slv(opcode_type, 16#07#),
      195 => to_slv(opcode_type, 16#02#),
      196 => to_slv(opcode_type, 16#0D#),
      197 => to_slv(opcode_type, 16#07#),
      198 => to_slv(opcode_type, 16#0D#),
      199 => to_slv(opcode_type, 16#11#),
      200 => to_slv(opcode_type, 16#09#),
      201 => to_slv(opcode_type, 16#01#),
      202 => to_slv(opcode_type, 16#08#),
      203 => to_slv(opcode_type, 16#10#),
      204 => to_slv(opcode_type, 16#0B#),
      205 => to_slv(opcode_type, 16#08#),
      206 => to_slv(opcode_type, 16#06#),
      207 => to_slv(opcode_type, 16#0C#),
      208 => to_slv(opcode_type, 16#0B#),
      209 => to_slv(opcode_type, 16#07#),
      210 => to_slv(opcode_type, 16#11#),
      211 => to_slv(opcode_type, 16#0D#),
      212 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#08#),
      225 => to_slv(opcode_type, 16#03#),
      226 => to_slv(opcode_type, 16#01#),
      227 => to_slv(opcode_type, 16#07#),
      228 => to_slv(opcode_type, 16#11#),
      229 => to_slv(opcode_type, 16#0D#),
      230 => to_slv(opcode_type, 16#07#),
      231 => to_slv(opcode_type, 16#08#),
      232 => to_slv(opcode_type, 16#08#),
      233 => to_slv(opcode_type, 16#0E#),
      234 => to_slv(opcode_type, 16#E0#),
      235 => to_slv(opcode_type, 16#06#),
      236 => to_slv(opcode_type, 16#0C#),
      237 => to_slv(opcode_type, 16#0A#),
      238 => to_slv(opcode_type, 16#09#),
      239 => to_slv(opcode_type, 16#08#),
      240 => to_slv(opcode_type, 16#0C#),
      241 => to_slv(opcode_type, 16#11#),
      242 => to_slv(opcode_type, 16#05#),
      243 => to_slv(opcode_type, 16#0C#),
      244 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#08#),
      257 => to_slv(opcode_type, 16#03#),
      258 => to_slv(opcode_type, 16#07#),
      259 => to_slv(opcode_type, 16#08#),
      260 => to_slv(opcode_type, 16#E8#),
      261 => to_slv(opcode_type, 16#0F#),
      262 => to_slv(opcode_type, 16#06#),
      263 => to_slv(opcode_type, 16#10#),
      264 => to_slv(opcode_type, 16#0B#),
      265 => to_slv(opcode_type, 16#07#),
      266 => to_slv(opcode_type, 16#09#),
      267 => to_slv(opcode_type, 16#03#),
      268 => to_slv(opcode_type, 16#0F#),
      269 => to_slv(opcode_type, 16#03#),
      270 => to_slv(opcode_type, 16#0D#),
      271 => to_slv(opcode_type, 16#08#),
      272 => to_slv(opcode_type, 16#09#),
      273 => to_slv(opcode_type, 16#10#),
      274 => to_slv(opcode_type, 16#0C#),
      275 => to_slv(opcode_type, 16#0B#),
      276 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#08#),
      289 => to_slv(opcode_type, 16#05#),
      290 => to_slv(opcode_type, 16#08#),
      291 => to_slv(opcode_type, 16#08#),
      292 => to_slv(opcode_type, 16#10#),
      293 => to_slv(opcode_type, 16#11#),
      294 => to_slv(opcode_type, 16#06#),
      295 => to_slv(opcode_type, 16#0F#),
      296 => to_slv(opcode_type, 16#11#),
      297 => to_slv(opcode_type, 16#09#),
      298 => to_slv(opcode_type, 16#07#),
      299 => to_slv(opcode_type, 16#04#),
      300 => to_slv(opcode_type, 16#0D#),
      301 => to_slv(opcode_type, 16#08#),
      302 => to_slv(opcode_type, 16#0A#),
      303 => to_slv(opcode_type, 16#D3#),
      304 => to_slv(opcode_type, 16#08#),
      305 => to_slv(opcode_type, 16#05#),
      306 => to_slv(opcode_type, 16#0F#),
      307 => to_slv(opcode_type, 16#0B#),
      308 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#09#),
      321 => to_slv(opcode_type, 16#04#),
      322 => to_slv(opcode_type, 16#09#),
      323 => to_slv(opcode_type, 16#07#),
      324 => to_slv(opcode_type, 16#0C#),
      325 => to_slv(opcode_type, 16#0D#),
      326 => to_slv(opcode_type, 16#06#),
      327 => to_slv(opcode_type, 16#0D#),
      328 => to_slv(opcode_type, 16#0D#),
      329 => to_slv(opcode_type, 16#09#),
      330 => to_slv(opcode_type, 16#02#),
      331 => to_slv(opcode_type, 16#06#),
      332 => to_slv(opcode_type, 16#0A#),
      333 => to_slv(opcode_type, 16#11#),
      334 => to_slv(opcode_type, 16#08#),
      335 => to_slv(opcode_type, 16#07#),
      336 => to_slv(opcode_type, 16#27#),
      337 => to_slv(opcode_type, 16#0B#),
      338 => to_slv(opcode_type, 16#02#),
      339 => to_slv(opcode_type, 16#0D#),
      340 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#07#),
      353 => to_slv(opcode_type, 16#07#),
      354 => to_slv(opcode_type, 16#08#),
      355 => to_slv(opcode_type, 16#08#),
      356 => to_slv(opcode_type, 16#10#),
      357 => to_slv(opcode_type, 16#B2#),
      358 => to_slv(opcode_type, 16#02#),
      359 => to_slv(opcode_type, 16#0D#),
      360 => to_slv(opcode_type, 16#05#),
      361 => to_slv(opcode_type, 16#05#),
      362 => to_slv(opcode_type, 16#10#),
      363 => to_slv(opcode_type, 16#08#),
      364 => to_slv(opcode_type, 16#09#),
      365 => to_slv(opcode_type, 16#01#),
      366 => to_slv(opcode_type, 16#0B#),
      367 => to_slv(opcode_type, 16#07#),
      368 => to_slv(opcode_type, 16#0F#),
      369 => to_slv(opcode_type, 16#0A#),
      370 => to_slv(opcode_type, 16#05#),
      371 => to_slv(opcode_type, 16#10#),
      372 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#07#),
      385 => to_slv(opcode_type, 16#08#),
      386 => to_slv(opcode_type, 16#04#),
      387 => to_slv(opcode_type, 16#08#),
      388 => to_slv(opcode_type, 16#0D#),
      389 => to_slv(opcode_type, 16#F7#),
      390 => to_slv(opcode_type, 16#04#),
      391 => to_slv(opcode_type, 16#02#),
      392 => to_slv(opcode_type, 16#10#),
      393 => to_slv(opcode_type, 16#08#),
      394 => to_slv(opcode_type, 16#06#),
      395 => to_slv(opcode_type, 16#06#),
      396 => to_slv(opcode_type, 16#0F#),
      397 => to_slv(opcode_type, 16#0F#),
      398 => to_slv(opcode_type, 16#06#),
      399 => to_slv(opcode_type, 16#10#),
      400 => to_slv(opcode_type, 16#6F#),
      401 => to_slv(opcode_type, 16#03#),
      402 => to_slv(opcode_type, 16#04#),
      403 => to_slv(opcode_type, 16#0B#),
      404 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#07#),
      417 => to_slv(opcode_type, 16#07#),
      418 => to_slv(opcode_type, 16#04#),
      419 => to_slv(opcode_type, 16#08#),
      420 => to_slv(opcode_type, 16#0D#),
      421 => to_slv(opcode_type, 16#10#),
      422 => to_slv(opcode_type, 16#09#),
      423 => to_slv(opcode_type, 16#02#),
      424 => to_slv(opcode_type, 16#11#),
      425 => to_slv(opcode_type, 16#04#),
      426 => to_slv(opcode_type, 16#10#),
      427 => to_slv(opcode_type, 16#07#),
      428 => to_slv(opcode_type, 16#04#),
      429 => to_slv(opcode_type, 16#03#),
      430 => to_slv(opcode_type, 16#0A#),
      431 => to_slv(opcode_type, 16#08#),
      432 => to_slv(opcode_type, 16#01#),
      433 => to_slv(opcode_type, 16#FD#),
      434 => to_slv(opcode_type, 16#01#),
      435 => to_slv(opcode_type, 16#0A#),
      436 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#07#),
      449 => to_slv(opcode_type, 16#01#),
      450 => to_slv(opcode_type, 16#06#),
      451 => to_slv(opcode_type, 16#09#),
      452 => to_slv(opcode_type, 16#8D#),
      453 => to_slv(opcode_type, 16#0D#),
      454 => to_slv(opcode_type, 16#09#),
      455 => to_slv(opcode_type, 16#0D#),
      456 => to_slv(opcode_type, 16#10#),
      457 => to_slv(opcode_type, 16#08#),
      458 => to_slv(opcode_type, 16#02#),
      459 => to_slv(opcode_type, 16#07#),
      460 => to_slv(opcode_type, 16#0A#),
      461 => to_slv(opcode_type, 16#11#),
      462 => to_slv(opcode_type, 16#08#),
      463 => to_slv(opcode_type, 16#08#),
      464 => to_slv(opcode_type, 16#0C#),
      465 => to_slv(opcode_type, 16#CB#),
      466 => to_slv(opcode_type, 16#03#),
      467 => to_slv(opcode_type, 16#29#),
      468 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#08#),
      481 => to_slv(opcode_type, 16#01#),
      482 => to_slv(opcode_type, 16#09#),
      483 => to_slv(opcode_type, 16#09#),
      484 => to_slv(opcode_type, 16#0C#),
      485 => to_slv(opcode_type, 16#EA#),
      486 => to_slv(opcode_type, 16#01#),
      487 => to_slv(opcode_type, 16#0C#),
      488 => to_slv(opcode_type, 16#09#),
      489 => to_slv(opcode_type, 16#09#),
      490 => to_slv(opcode_type, 16#06#),
      491 => to_slv(opcode_type, 16#11#),
      492 => to_slv(opcode_type, 16#10#),
      493 => to_slv(opcode_type, 16#08#),
      494 => to_slv(opcode_type, 16#10#),
      495 => to_slv(opcode_type, 16#0D#),
      496 => to_slv(opcode_type, 16#08#),
      497 => to_slv(opcode_type, 16#05#),
      498 => to_slv(opcode_type, 16#10#),
      499 => to_slv(opcode_type, 16#0F#),
      500 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#06#),
      513 => to_slv(opcode_type, 16#02#),
      514 => to_slv(opcode_type, 16#08#),
      515 => to_slv(opcode_type, 16#04#),
      516 => to_slv(opcode_type, 16#11#),
      517 => to_slv(opcode_type, 16#01#),
      518 => to_slv(opcode_type, 16#0C#),
      519 => to_slv(opcode_type, 16#07#),
      520 => to_slv(opcode_type, 16#07#),
      521 => to_slv(opcode_type, 16#02#),
      522 => to_slv(opcode_type, 16#0F#),
      523 => to_slv(opcode_type, 16#01#),
      524 => to_slv(opcode_type, 16#0C#),
      525 => to_slv(opcode_type, 16#07#),
      526 => to_slv(opcode_type, 16#06#),
      527 => to_slv(opcode_type, 16#0A#),
      528 => to_slv(opcode_type, 16#0D#),
      529 => to_slv(opcode_type, 16#07#),
      530 => to_slv(opcode_type, 16#9B#),
      531 => to_slv(opcode_type, 16#0B#),
      532 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#09#),
      545 => to_slv(opcode_type, 16#07#),
      546 => to_slv(opcode_type, 16#07#),
      547 => to_slv(opcode_type, 16#01#),
      548 => to_slv(opcode_type, 16#0C#),
      549 => to_slv(opcode_type, 16#06#),
      550 => to_slv(opcode_type, 16#11#),
      551 => to_slv(opcode_type, 16#1E#),
      552 => to_slv(opcode_type, 16#02#),
      553 => to_slv(opcode_type, 16#07#),
      554 => to_slv(opcode_type, 16#0F#),
      555 => to_slv(opcode_type, 16#0A#),
      556 => to_slv(opcode_type, 16#09#),
      557 => to_slv(opcode_type, 16#04#),
      558 => to_slv(opcode_type, 16#07#),
      559 => to_slv(opcode_type, 16#0D#),
      560 => to_slv(opcode_type, 16#11#),
      561 => to_slv(opcode_type, 16#04#),
      562 => to_slv(opcode_type, 16#03#),
      563 => to_slv(opcode_type, 16#11#),
      564 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#08#),
      577 => to_slv(opcode_type, 16#03#),
      578 => to_slv(opcode_type, 16#03#),
      579 => to_slv(opcode_type, 16#07#),
      580 => to_slv(opcode_type, 16#0A#),
      581 => to_slv(opcode_type, 16#0B#),
      582 => to_slv(opcode_type, 16#07#),
      583 => to_slv(opcode_type, 16#07#),
      584 => to_slv(opcode_type, 16#08#),
      585 => to_slv(opcode_type, 16#0B#),
      586 => to_slv(opcode_type, 16#0F#),
      587 => to_slv(opcode_type, 16#03#),
      588 => to_slv(opcode_type, 16#11#),
      589 => to_slv(opcode_type, 16#08#),
      590 => to_slv(opcode_type, 16#09#),
      591 => to_slv(opcode_type, 16#11#),
      592 => to_slv(opcode_type, 16#0D#),
      593 => to_slv(opcode_type, 16#09#),
      594 => to_slv(opcode_type, 16#11#),
      595 => to_slv(opcode_type, 16#0A#),
      596 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#06#),
      609 => to_slv(opcode_type, 16#05#),
      610 => to_slv(opcode_type, 16#07#),
      611 => to_slv(opcode_type, 16#04#),
      612 => to_slv(opcode_type, 16#0B#),
      613 => to_slv(opcode_type, 16#05#),
      614 => to_slv(opcode_type, 16#0E#),
      615 => to_slv(opcode_type, 16#07#),
      616 => to_slv(opcode_type, 16#06#),
      617 => to_slv(opcode_type, 16#01#),
      618 => to_slv(opcode_type, 16#0F#),
      619 => to_slv(opcode_type, 16#05#),
      620 => to_slv(opcode_type, 16#0F#),
      621 => to_slv(opcode_type, 16#09#),
      622 => to_slv(opcode_type, 16#07#),
      623 => to_slv(opcode_type, 16#0A#),
      624 => to_slv(opcode_type, 16#11#),
      625 => to_slv(opcode_type, 16#08#),
      626 => to_slv(opcode_type, 16#10#),
      627 => to_slv(opcode_type, 16#0F#),
      628 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#08#),
      641 => to_slv(opcode_type, 16#09#),
      642 => to_slv(opcode_type, 16#01#),
      643 => to_slv(opcode_type, 16#06#),
      644 => to_slv(opcode_type, 16#0D#),
      645 => to_slv(opcode_type, 16#0B#),
      646 => to_slv(opcode_type, 16#04#),
      647 => to_slv(opcode_type, 16#02#),
      648 => to_slv(opcode_type, 16#11#),
      649 => to_slv(opcode_type, 16#07#),
      650 => to_slv(opcode_type, 16#09#),
      651 => to_slv(opcode_type, 16#08#),
      652 => to_slv(opcode_type, 16#0A#),
      653 => to_slv(opcode_type, 16#0A#),
      654 => to_slv(opcode_type, 16#06#),
      655 => to_slv(opcode_type, 16#0C#),
      656 => to_slv(opcode_type, 16#0A#),
      657 => to_slv(opcode_type, 16#06#),
      658 => to_slv(opcode_type, 16#0B#),
      659 => to_slv(opcode_type, 16#0E#),
      660 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#06#),
      673 => to_slv(opcode_type, 16#04#),
      674 => to_slv(opcode_type, 16#01#),
      675 => to_slv(opcode_type, 16#04#),
      676 => to_slv(opcode_type, 16#0D#),
      677 => to_slv(opcode_type, 16#08#),
      678 => to_slv(opcode_type, 16#07#),
      679 => to_slv(opcode_type, 16#07#),
      680 => to_slv(opcode_type, 16#11#),
      681 => to_slv(opcode_type, 16#0E#),
      682 => to_slv(opcode_type, 16#08#),
      683 => to_slv(opcode_type, 16#0D#),
      684 => to_slv(opcode_type, 16#10#),
      685 => to_slv(opcode_type, 16#07#),
      686 => to_slv(opcode_type, 16#07#),
      687 => to_slv(opcode_type, 16#0F#),
      688 => to_slv(opcode_type, 16#0B#),
      689 => to_slv(opcode_type, 16#08#),
      690 => to_slv(opcode_type, 16#0B#),
      691 => to_slv(opcode_type, 16#0D#),
      692 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#06#),
      705 => to_slv(opcode_type, 16#09#),
      706 => to_slv(opcode_type, 16#03#),
      707 => to_slv(opcode_type, 16#08#),
      708 => to_slv(opcode_type, 16#10#),
      709 => to_slv(opcode_type, 16#10#),
      710 => to_slv(opcode_type, 16#05#),
      711 => to_slv(opcode_type, 16#08#),
      712 => to_slv(opcode_type, 16#75#),
      713 => to_slv(opcode_type, 16#0A#),
      714 => to_slv(opcode_type, 16#06#),
      715 => to_slv(opcode_type, 16#07#),
      716 => to_slv(opcode_type, 16#06#),
      717 => to_slv(opcode_type, 16#2A#),
      718 => to_slv(opcode_type, 16#0C#),
      719 => to_slv(opcode_type, 16#01#),
      720 => to_slv(opcode_type, 16#0A#),
      721 => to_slv(opcode_type, 16#07#),
      722 => to_slv(opcode_type, 16#11#),
      723 => to_slv(opcode_type, 16#0E#),
      724 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#09#),
      737 => to_slv(opcode_type, 16#07#),
      738 => to_slv(opcode_type, 16#07#),
      739 => to_slv(opcode_type, 16#01#),
      740 => to_slv(opcode_type, 16#0A#),
      741 => to_slv(opcode_type, 16#04#),
      742 => to_slv(opcode_type, 16#0E#),
      743 => to_slv(opcode_type, 16#08#),
      744 => to_slv(opcode_type, 16#05#),
      745 => to_slv(opcode_type, 16#0E#),
      746 => to_slv(opcode_type, 16#09#),
      747 => to_slv(opcode_type, 16#0A#),
      748 => to_slv(opcode_type, 16#0C#),
      749 => to_slv(opcode_type, 16#09#),
      750 => to_slv(opcode_type, 16#04#),
      751 => to_slv(opcode_type, 16#03#),
      752 => to_slv(opcode_type, 16#0E#),
      753 => to_slv(opcode_type, 16#09#),
      754 => to_slv(opcode_type, 16#11#),
      755 => to_slv(opcode_type, 16#0F#),
      756 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#07#),
      769 => to_slv(opcode_type, 16#04#),
      770 => to_slv(opcode_type, 16#02#),
      771 => to_slv(opcode_type, 16#05#),
      772 => to_slv(opcode_type, 16#0D#),
      773 => to_slv(opcode_type, 16#07#),
      774 => to_slv(opcode_type, 16#08#),
      775 => to_slv(opcode_type, 16#07#),
      776 => to_slv(opcode_type, 16#0F#),
      777 => to_slv(opcode_type, 16#0E#),
      778 => to_slv(opcode_type, 16#07#),
      779 => to_slv(opcode_type, 16#0F#),
      780 => to_slv(opcode_type, 16#0C#),
      781 => to_slv(opcode_type, 16#07#),
      782 => to_slv(opcode_type, 16#08#),
      783 => to_slv(opcode_type, 16#0B#),
      784 => to_slv(opcode_type, 16#10#),
      785 => to_slv(opcode_type, 16#06#),
      786 => to_slv(opcode_type, 16#10#),
      787 => to_slv(opcode_type, 16#0B#),
      788 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#09#),
      801 => to_slv(opcode_type, 16#04#),
      802 => to_slv(opcode_type, 16#01#),
      803 => to_slv(opcode_type, 16#02#),
      804 => to_slv(opcode_type, 16#10#),
      805 => to_slv(opcode_type, 16#06#),
      806 => to_slv(opcode_type, 16#09#),
      807 => to_slv(opcode_type, 16#07#),
      808 => to_slv(opcode_type, 16#0C#),
      809 => to_slv(opcode_type, 16#0B#),
      810 => to_slv(opcode_type, 16#07#),
      811 => to_slv(opcode_type, 16#0B#),
      812 => to_slv(opcode_type, 16#0A#),
      813 => to_slv(opcode_type, 16#09#),
      814 => to_slv(opcode_type, 16#09#),
      815 => to_slv(opcode_type, 16#0B#),
      816 => to_slv(opcode_type, 16#0C#),
      817 => to_slv(opcode_type, 16#07#),
      818 => to_slv(opcode_type, 16#0C#),
      819 => to_slv(opcode_type, 16#0A#),
      820 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#06#),
      833 => to_slv(opcode_type, 16#06#),
      834 => to_slv(opcode_type, 16#07#),
      835 => to_slv(opcode_type, 16#05#),
      836 => to_slv(opcode_type, 16#0F#),
      837 => to_slv(opcode_type, 16#09#),
      838 => to_slv(opcode_type, 16#0E#),
      839 => to_slv(opcode_type, 16#11#),
      840 => to_slv(opcode_type, 16#08#),
      841 => to_slv(opcode_type, 16#06#),
      842 => to_slv(opcode_type, 16#0F#),
      843 => to_slv(opcode_type, 16#0F#),
      844 => to_slv(opcode_type, 16#07#),
      845 => to_slv(opcode_type, 16#0F#),
      846 => to_slv(opcode_type, 16#0B#),
      847 => to_slv(opcode_type, 16#03#),
      848 => to_slv(opcode_type, 16#07#),
      849 => to_slv(opcode_type, 16#05#),
      850 => to_slv(opcode_type, 16#0C#),
      851 => to_slv(opcode_type, 16#10#),
      852 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#06#),
      865 => to_slv(opcode_type, 16#03#),
      866 => to_slv(opcode_type, 16#04#),
      867 => to_slv(opcode_type, 16#09#),
      868 => to_slv(opcode_type, 16#11#),
      869 => to_slv(opcode_type, 16#0C#),
      870 => to_slv(opcode_type, 16#08#),
      871 => to_slv(opcode_type, 16#06#),
      872 => to_slv(opcode_type, 16#06#),
      873 => to_slv(opcode_type, 16#0D#),
      874 => to_slv(opcode_type, 16#DC#),
      875 => to_slv(opcode_type, 16#07#),
      876 => to_slv(opcode_type, 16#0A#),
      877 => to_slv(opcode_type, 16#0B#),
      878 => to_slv(opcode_type, 16#07#),
      879 => to_slv(opcode_type, 16#02#),
      880 => to_slv(opcode_type, 16#10#),
      881 => to_slv(opcode_type, 16#06#),
      882 => to_slv(opcode_type, 16#11#),
      883 => to_slv(opcode_type, 16#0E#),
      884 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#09#),
      897 => to_slv(opcode_type, 16#08#),
      898 => to_slv(opcode_type, 16#03#),
      899 => to_slv(opcode_type, 16#09#),
      900 => to_slv(opcode_type, 16#0A#),
      901 => to_slv(opcode_type, 16#11#),
      902 => to_slv(opcode_type, 16#07#),
      903 => to_slv(opcode_type, 16#04#),
      904 => to_slv(opcode_type, 16#11#),
      905 => to_slv(opcode_type, 16#04#),
      906 => to_slv(opcode_type, 16#11#),
      907 => to_slv(opcode_type, 16#08#),
      908 => to_slv(opcode_type, 16#04#),
      909 => to_slv(opcode_type, 16#04#),
      910 => to_slv(opcode_type, 16#0F#),
      911 => to_slv(opcode_type, 16#07#),
      912 => to_slv(opcode_type, 16#05#),
      913 => to_slv(opcode_type, 16#C0#),
      914 => to_slv(opcode_type, 16#02#),
      915 => to_slv(opcode_type, 16#0B#),
      916 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#09#),
      929 => to_slv(opcode_type, 16#04#),
      930 => to_slv(opcode_type, 16#04#),
      931 => to_slv(opcode_type, 16#08#),
      932 => to_slv(opcode_type, 16#0D#),
      933 => to_slv(opcode_type, 16#10#),
      934 => to_slv(opcode_type, 16#07#),
      935 => to_slv(opcode_type, 16#07#),
      936 => to_slv(opcode_type, 16#06#),
      937 => to_slv(opcode_type, 16#0E#),
      938 => to_slv(opcode_type, 16#0D#),
      939 => to_slv(opcode_type, 16#07#),
      940 => to_slv(opcode_type, 16#8C#),
      941 => to_slv(opcode_type, 16#0A#),
      942 => to_slv(opcode_type, 16#08#),
      943 => to_slv(opcode_type, 16#01#),
      944 => to_slv(opcode_type, 16#14#),
      945 => to_slv(opcode_type, 16#08#),
      946 => to_slv(opcode_type, 16#0A#),
      947 => to_slv(opcode_type, 16#11#),
      948 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#09#),
      961 => to_slv(opcode_type, 16#07#),
      962 => to_slv(opcode_type, 16#04#),
      963 => to_slv(opcode_type, 16#04#),
      964 => to_slv(opcode_type, 16#11#),
      965 => to_slv(opcode_type, 16#07#),
      966 => to_slv(opcode_type, 16#03#),
      967 => to_slv(opcode_type, 16#0B#),
      968 => to_slv(opcode_type, 16#05#),
      969 => to_slv(opcode_type, 16#0C#),
      970 => to_slv(opcode_type, 16#07#),
      971 => to_slv(opcode_type, 16#02#),
      972 => to_slv(opcode_type, 16#06#),
      973 => to_slv(opcode_type, 16#0A#),
      974 => to_slv(opcode_type, 16#0B#),
      975 => to_slv(opcode_type, 16#07#),
      976 => to_slv(opcode_type, 16#07#),
      977 => to_slv(opcode_type, 16#0A#),
      978 => to_slv(opcode_type, 16#0E#),
      979 => to_slv(opcode_type, 16#0A#),
      980 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#08#),
      993 => to_slv(opcode_type, 16#09#),
      994 => to_slv(opcode_type, 16#07#),
      995 => to_slv(opcode_type, 16#02#),
      996 => to_slv(opcode_type, 16#0A#),
      997 => to_slv(opcode_type, 16#09#),
      998 => to_slv(opcode_type, 16#10#),
      999 => to_slv(opcode_type, 16#10#),
      1000 => to_slv(opcode_type, 16#09#),
      1001 => to_slv(opcode_type, 16#08#),
      1002 => to_slv(opcode_type, 16#0D#),
      1003 => to_slv(opcode_type, 16#0D#),
      1004 => to_slv(opcode_type, 16#02#),
      1005 => to_slv(opcode_type, 16#10#),
      1006 => to_slv(opcode_type, 16#07#),
      1007 => to_slv(opcode_type, 16#05#),
      1008 => to_slv(opcode_type, 16#06#),
      1009 => to_slv(opcode_type, 16#0C#),
      1010 => to_slv(opcode_type, 16#0E#),
      1011 => to_slv(opcode_type, 16#10#),
      1012 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#07#),
      1025 => to_slv(opcode_type, 16#05#),
      1026 => to_slv(opcode_type, 16#08#),
      1027 => to_slv(opcode_type, 16#03#),
      1028 => to_slv(opcode_type, 16#0A#),
      1029 => to_slv(opcode_type, 16#01#),
      1030 => to_slv(opcode_type, 16#0C#),
      1031 => to_slv(opcode_type, 16#07#),
      1032 => to_slv(opcode_type, 16#09#),
      1033 => to_slv(opcode_type, 16#03#),
      1034 => to_slv(opcode_type, 16#0D#),
      1035 => to_slv(opcode_type, 16#07#),
      1036 => to_slv(opcode_type, 16#0A#),
      1037 => to_slv(opcode_type, 16#10#),
      1038 => to_slv(opcode_type, 16#07#),
      1039 => to_slv(opcode_type, 16#09#),
      1040 => to_slv(opcode_type, 16#0D#),
      1041 => to_slv(opcode_type, 16#0E#),
      1042 => to_slv(opcode_type, 16#02#),
      1043 => to_slv(opcode_type, 16#0B#),
      1044 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#07#),
      1057 => to_slv(opcode_type, 16#01#),
      1058 => to_slv(opcode_type, 16#01#),
      1059 => to_slv(opcode_type, 16#07#),
      1060 => to_slv(opcode_type, 16#0A#),
      1061 => to_slv(opcode_type, 16#98#),
      1062 => to_slv(opcode_type, 16#08#),
      1063 => to_slv(opcode_type, 16#08#),
      1064 => to_slv(opcode_type, 16#02#),
      1065 => to_slv(opcode_type, 16#0D#),
      1066 => to_slv(opcode_type, 16#09#),
      1067 => to_slv(opcode_type, 16#0B#),
      1068 => to_slv(opcode_type, 16#10#),
      1069 => to_slv(opcode_type, 16#06#),
      1070 => to_slv(opcode_type, 16#07#),
      1071 => to_slv(opcode_type, 16#0E#),
      1072 => to_slv(opcode_type, 16#0D#),
      1073 => to_slv(opcode_type, 16#06#),
      1074 => to_slv(opcode_type, 16#0A#),
      1075 => to_slv(opcode_type, 16#0E#),
      1076 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#06#),
      1089 => to_slv(opcode_type, 16#03#),
      1090 => to_slv(opcode_type, 16#07#),
      1091 => to_slv(opcode_type, 16#08#),
      1092 => to_slv(opcode_type, 16#10#),
      1093 => to_slv(opcode_type, 16#0E#),
      1094 => to_slv(opcode_type, 16#04#),
      1095 => to_slv(opcode_type, 16#0D#),
      1096 => to_slv(opcode_type, 16#08#),
      1097 => to_slv(opcode_type, 16#01#),
      1098 => to_slv(opcode_type, 16#07#),
      1099 => to_slv(opcode_type, 16#0D#),
      1100 => to_slv(opcode_type, 16#0C#),
      1101 => to_slv(opcode_type, 16#07#),
      1102 => to_slv(opcode_type, 16#07#),
      1103 => to_slv(opcode_type, 16#10#),
      1104 => to_slv(opcode_type, 16#0F#),
      1105 => to_slv(opcode_type, 16#06#),
      1106 => to_slv(opcode_type, 16#0F#),
      1107 => to_slv(opcode_type, 16#0C#),
      1108 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#07#),
      1121 => to_slv(opcode_type, 16#03#),
      1122 => to_slv(opcode_type, 16#08#),
      1123 => to_slv(opcode_type, 16#08#),
      1124 => to_slv(opcode_type, 16#10#),
      1125 => to_slv(opcode_type, 16#0F#),
      1126 => to_slv(opcode_type, 16#06#),
      1127 => to_slv(opcode_type, 16#0C#),
      1128 => to_slv(opcode_type, 16#0C#),
      1129 => to_slv(opcode_type, 16#08#),
      1130 => to_slv(opcode_type, 16#09#),
      1131 => to_slv(opcode_type, 16#01#),
      1132 => to_slv(opcode_type, 16#0D#),
      1133 => to_slv(opcode_type, 16#02#),
      1134 => to_slv(opcode_type, 16#0D#),
      1135 => to_slv(opcode_type, 16#09#),
      1136 => to_slv(opcode_type, 16#09#),
      1137 => to_slv(opcode_type, 16#0A#),
      1138 => to_slv(opcode_type, 16#0C#),
      1139 => to_slv(opcode_type, 16#0C#),
      1140 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#07#),
      1153 => to_slv(opcode_type, 16#08#),
      1154 => to_slv(opcode_type, 16#06#),
      1155 => to_slv(opcode_type, 16#06#),
      1156 => to_slv(opcode_type, 16#0F#),
      1157 => to_slv(opcode_type, 16#0E#),
      1158 => to_slv(opcode_type, 16#03#),
      1159 => to_slv(opcode_type, 16#0B#),
      1160 => to_slv(opcode_type, 16#02#),
      1161 => to_slv(opcode_type, 16#02#),
      1162 => to_slv(opcode_type, 16#0F#),
      1163 => to_slv(opcode_type, 16#07#),
      1164 => to_slv(opcode_type, 16#06#),
      1165 => to_slv(opcode_type, 16#06#),
      1166 => to_slv(opcode_type, 16#10#),
      1167 => to_slv(opcode_type, 16#0D#),
      1168 => to_slv(opcode_type, 16#04#),
      1169 => to_slv(opcode_type, 16#0A#),
      1170 => to_slv(opcode_type, 16#04#),
      1171 => to_slv(opcode_type, 16#0D#),
      1172 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#06#),
      1185 => to_slv(opcode_type, 16#01#),
      1186 => to_slv(opcode_type, 16#09#),
      1187 => to_slv(opcode_type, 16#09#),
      1188 => to_slv(opcode_type, 16#E7#),
      1189 => to_slv(opcode_type, 16#0A#),
      1190 => to_slv(opcode_type, 16#06#),
      1191 => to_slv(opcode_type, 16#10#),
      1192 => to_slv(opcode_type, 16#0F#),
      1193 => to_slv(opcode_type, 16#07#),
      1194 => to_slv(opcode_type, 16#06#),
      1195 => to_slv(opcode_type, 16#01#),
      1196 => to_slv(opcode_type, 16#0B#),
      1197 => to_slv(opcode_type, 16#09#),
      1198 => to_slv(opcode_type, 16#10#),
      1199 => to_slv(opcode_type, 16#14#),
      1200 => to_slv(opcode_type, 16#01#),
      1201 => to_slv(opcode_type, 16#09#),
      1202 => to_slv(opcode_type, 16#0B#),
      1203 => to_slv(opcode_type, 16#0A#),
      1204 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#08#),
      1217 => to_slv(opcode_type, 16#02#),
      1218 => to_slv(opcode_type, 16#06#),
      1219 => to_slv(opcode_type, 16#08#),
      1220 => to_slv(opcode_type, 16#11#),
      1221 => to_slv(opcode_type, 16#0F#),
      1222 => to_slv(opcode_type, 16#03#),
      1223 => to_slv(opcode_type, 16#0D#),
      1224 => to_slv(opcode_type, 16#08#),
      1225 => to_slv(opcode_type, 16#09#),
      1226 => to_slv(opcode_type, 16#02#),
      1227 => to_slv(opcode_type, 16#0F#),
      1228 => to_slv(opcode_type, 16#04#),
      1229 => to_slv(opcode_type, 16#10#),
      1230 => to_slv(opcode_type, 16#07#),
      1231 => to_slv(opcode_type, 16#04#),
      1232 => to_slv(opcode_type, 16#0C#),
      1233 => to_slv(opcode_type, 16#06#),
      1234 => to_slv(opcode_type, 16#0F#),
      1235 => to_slv(opcode_type, 16#0E#),
      1236 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#09#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#04#),
      1251 => to_slv(opcode_type, 16#05#),
      1252 => to_slv(opcode_type, 16#11#),
      1253 => to_slv(opcode_type, 16#02#),
      1254 => to_slv(opcode_type, 16#03#),
      1255 => to_slv(opcode_type, 16#0C#),
      1256 => to_slv(opcode_type, 16#09#),
      1257 => to_slv(opcode_type, 16#06#),
      1258 => to_slv(opcode_type, 16#09#),
      1259 => to_slv(opcode_type, 16#11#),
      1260 => to_slv(opcode_type, 16#0E#),
      1261 => to_slv(opcode_type, 16#04#),
      1262 => to_slv(opcode_type, 16#0B#),
      1263 => to_slv(opcode_type, 16#06#),
      1264 => to_slv(opcode_type, 16#06#),
      1265 => to_slv(opcode_type, 16#10#),
      1266 => to_slv(opcode_type, 16#11#),
      1267 => to_slv(opcode_type, 16#0C#),
      1268 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#08#),
      1281 => to_slv(opcode_type, 16#02#),
      1282 => to_slv(opcode_type, 16#09#),
      1283 => to_slv(opcode_type, 16#06#),
      1284 => to_slv(opcode_type, 16#11#),
      1285 => to_slv(opcode_type, 16#0D#),
      1286 => to_slv(opcode_type, 16#05#),
      1287 => to_slv(opcode_type, 16#0A#),
      1288 => to_slv(opcode_type, 16#06#),
      1289 => to_slv(opcode_type, 16#05#),
      1290 => to_slv(opcode_type, 16#08#),
      1291 => to_slv(opcode_type, 16#10#),
      1292 => to_slv(opcode_type, 16#B3#),
      1293 => to_slv(opcode_type, 16#07#),
      1294 => to_slv(opcode_type, 16#07#),
      1295 => to_slv(opcode_type, 16#E5#),
      1296 => to_slv(opcode_type, 16#F7#),
      1297 => to_slv(opcode_type, 16#07#),
      1298 => to_slv(opcode_type, 16#0A#),
      1299 => to_slv(opcode_type, 16#0E#),
      1300 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#09#),
      1313 => to_slv(opcode_type, 16#01#),
      1314 => to_slv(opcode_type, 16#08#),
      1315 => to_slv(opcode_type, 16#09#),
      1316 => to_slv(opcode_type, 16#0D#),
      1317 => to_slv(opcode_type, 16#0D#),
      1318 => to_slv(opcode_type, 16#02#),
      1319 => to_slv(opcode_type, 16#0E#),
      1320 => to_slv(opcode_type, 16#08#),
      1321 => to_slv(opcode_type, 16#07#),
      1322 => to_slv(opcode_type, 16#05#),
      1323 => to_slv(opcode_type, 16#0E#),
      1324 => to_slv(opcode_type, 16#01#),
      1325 => to_slv(opcode_type, 16#0D#),
      1326 => to_slv(opcode_type, 16#07#),
      1327 => to_slv(opcode_type, 16#05#),
      1328 => to_slv(opcode_type, 16#0B#),
      1329 => to_slv(opcode_type, 16#07#),
      1330 => to_slv(opcode_type, 16#0C#),
      1331 => to_slv(opcode_type, 16#11#),
      1332 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#08#),
      1345 => to_slv(opcode_type, 16#06#),
      1346 => to_slv(opcode_type, 16#08#),
      1347 => to_slv(opcode_type, 16#02#),
      1348 => to_slv(opcode_type, 16#0E#),
      1349 => to_slv(opcode_type, 16#08#),
      1350 => to_slv(opcode_type, 16#C6#),
      1351 => to_slv(opcode_type, 16#0B#),
      1352 => to_slv(opcode_type, 16#07#),
      1353 => to_slv(opcode_type, 16#07#),
      1354 => to_slv(opcode_type, 16#0B#),
      1355 => to_slv(opcode_type, 16#0C#),
      1356 => to_slv(opcode_type, 16#09#),
      1357 => to_slv(opcode_type, 16#0F#),
      1358 => to_slv(opcode_type, 16#10#),
      1359 => to_slv(opcode_type, 16#06#),
      1360 => to_slv(opcode_type, 16#02#),
      1361 => to_slv(opcode_type, 16#05#),
      1362 => to_slv(opcode_type, 16#0C#),
      1363 => to_slv(opcode_type, 16#0D#),
      1364 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#09#),
      1377 => to_slv(opcode_type, 16#09#),
      1378 => to_slv(opcode_type, 16#06#),
      1379 => to_slv(opcode_type, 16#07#),
      1380 => to_slv(opcode_type, 16#0B#),
      1381 => to_slv(opcode_type, 16#0E#),
      1382 => to_slv(opcode_type, 16#08#),
      1383 => to_slv(opcode_type, 16#0B#),
      1384 => to_slv(opcode_type, 16#0B#),
      1385 => to_slv(opcode_type, 16#07#),
      1386 => to_slv(opcode_type, 16#09#),
      1387 => to_slv(opcode_type, 16#0A#),
      1388 => to_slv(opcode_type, 16#0B#),
      1389 => to_slv(opcode_type, 16#01#),
      1390 => to_slv(opcode_type, 16#77#),
      1391 => to_slv(opcode_type, 16#09#),
      1392 => to_slv(opcode_type, 16#02#),
      1393 => to_slv(opcode_type, 16#03#),
      1394 => to_slv(opcode_type, 16#11#),
      1395 => to_slv(opcode_type, 16#50#),
      1396 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#09#),
      1409 => to_slv(opcode_type, 16#09#),
      1410 => to_slv(opcode_type, 16#01#),
      1411 => to_slv(opcode_type, 16#09#),
      1412 => to_slv(opcode_type, 16#FF#),
      1413 => to_slv(opcode_type, 16#0D#),
      1414 => to_slv(opcode_type, 16#09#),
      1415 => to_slv(opcode_type, 16#08#),
      1416 => to_slv(opcode_type, 16#0F#),
      1417 => to_slv(opcode_type, 16#0F#),
      1418 => to_slv(opcode_type, 16#09#),
      1419 => to_slv(opcode_type, 16#0E#),
      1420 => to_slv(opcode_type, 16#11#),
      1421 => to_slv(opcode_type, 16#07#),
      1422 => to_slv(opcode_type, 16#05#),
      1423 => to_slv(opcode_type, 16#09#),
      1424 => to_slv(opcode_type, 16#11#),
      1425 => to_slv(opcode_type, 16#0A#),
      1426 => to_slv(opcode_type, 16#03#),
      1427 => to_slv(opcode_type, 16#0D#),
      1428 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#07#),
      1441 => to_slv(opcode_type, 16#05#),
      1442 => to_slv(opcode_type, 16#06#),
      1443 => to_slv(opcode_type, 16#03#),
      1444 => to_slv(opcode_type, 16#0B#),
      1445 => to_slv(opcode_type, 16#08#),
      1446 => to_slv(opcode_type, 16#0C#),
      1447 => to_slv(opcode_type, 16#0B#),
      1448 => to_slv(opcode_type, 16#08#),
      1449 => to_slv(opcode_type, 16#01#),
      1450 => to_slv(opcode_type, 16#08#),
      1451 => to_slv(opcode_type, 16#0F#),
      1452 => to_slv(opcode_type, 16#11#),
      1453 => to_slv(opcode_type, 16#06#),
      1454 => to_slv(opcode_type, 16#08#),
      1455 => to_slv(opcode_type, 16#0E#),
      1456 => to_slv(opcode_type, 16#0C#),
      1457 => to_slv(opcode_type, 16#06#),
      1458 => to_slv(opcode_type, 16#0F#),
      1459 => to_slv(opcode_type, 16#0E#),
      1460 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#09#),
      1473 => to_slv(opcode_type, 16#08#),
      1474 => to_slv(opcode_type, 16#08#),
      1475 => to_slv(opcode_type, 16#09#),
      1476 => to_slv(opcode_type, 16#0E#),
      1477 => to_slv(opcode_type, 16#0C#),
      1478 => to_slv(opcode_type, 16#01#),
      1479 => to_slv(opcode_type, 16#0A#),
      1480 => to_slv(opcode_type, 16#05#),
      1481 => to_slv(opcode_type, 16#04#),
      1482 => to_slv(opcode_type, 16#0F#),
      1483 => to_slv(opcode_type, 16#08#),
      1484 => to_slv(opcode_type, 16#04#),
      1485 => to_slv(opcode_type, 16#04#),
      1486 => to_slv(opcode_type, 16#0F#),
      1487 => to_slv(opcode_type, 16#07#),
      1488 => to_slv(opcode_type, 16#03#),
      1489 => to_slv(opcode_type, 16#0D#),
      1490 => to_slv(opcode_type, 16#05#),
      1491 => to_slv(opcode_type, 16#0D#),
      1492 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#09#),
      1505 => to_slv(opcode_type, 16#07#),
      1506 => to_slv(opcode_type, 16#05#),
      1507 => to_slv(opcode_type, 16#08#),
      1508 => to_slv(opcode_type, 16#10#),
      1509 => to_slv(opcode_type, 16#0F#),
      1510 => to_slv(opcode_type, 16#05#),
      1511 => to_slv(opcode_type, 16#04#),
      1512 => to_slv(opcode_type, 16#0F#),
      1513 => to_slv(opcode_type, 16#07#),
      1514 => to_slv(opcode_type, 16#07#),
      1515 => to_slv(opcode_type, 16#03#),
      1516 => to_slv(opcode_type, 16#0B#),
      1517 => to_slv(opcode_type, 16#05#),
      1518 => to_slv(opcode_type, 16#0C#),
      1519 => to_slv(opcode_type, 16#07#),
      1520 => to_slv(opcode_type, 16#09#),
      1521 => to_slv(opcode_type, 16#0C#),
      1522 => to_slv(opcode_type, 16#0C#),
      1523 => to_slv(opcode_type, 16#1D#),
      1524 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#06#),
      1537 => to_slv(opcode_type, 16#09#),
      1538 => to_slv(opcode_type, 16#08#),
      1539 => to_slv(opcode_type, 16#05#),
      1540 => to_slv(opcode_type, 16#0B#),
      1541 => to_slv(opcode_type, 16#05#),
      1542 => to_slv(opcode_type, 16#0C#),
      1543 => to_slv(opcode_type, 16#08#),
      1544 => to_slv(opcode_type, 16#08#),
      1545 => to_slv(opcode_type, 16#0F#),
      1546 => to_slv(opcode_type, 16#0B#),
      1547 => to_slv(opcode_type, 16#05#),
      1548 => to_slv(opcode_type, 16#10#),
      1549 => to_slv(opcode_type, 16#04#),
      1550 => to_slv(opcode_type, 16#07#),
      1551 => to_slv(opcode_type, 16#02#),
      1552 => to_slv(opcode_type, 16#6C#),
      1553 => to_slv(opcode_type, 16#07#),
      1554 => to_slv(opcode_type, 16#0F#),
      1555 => to_slv(opcode_type, 16#0C#),
      1556 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#08#),
      1569 => to_slv(opcode_type, 16#03#),
      1570 => to_slv(opcode_type, 16#03#),
      1571 => to_slv(opcode_type, 16#05#),
      1572 => to_slv(opcode_type, 16#0E#),
      1573 => to_slv(opcode_type, 16#07#),
      1574 => to_slv(opcode_type, 16#07#),
      1575 => to_slv(opcode_type, 16#09#),
      1576 => to_slv(opcode_type, 16#0F#),
      1577 => to_slv(opcode_type, 16#0A#),
      1578 => to_slv(opcode_type, 16#06#),
      1579 => to_slv(opcode_type, 16#0B#),
      1580 => to_slv(opcode_type, 16#10#),
      1581 => to_slv(opcode_type, 16#09#),
      1582 => to_slv(opcode_type, 16#07#),
      1583 => to_slv(opcode_type, 16#0D#),
      1584 => to_slv(opcode_type, 16#0E#),
      1585 => to_slv(opcode_type, 16#06#),
      1586 => to_slv(opcode_type, 16#0E#),
      1587 => to_slv(opcode_type, 16#0F#),
      1588 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#07#),
      1601 => to_slv(opcode_type, 16#04#),
      1602 => to_slv(opcode_type, 16#06#),
      1603 => to_slv(opcode_type, 16#04#),
      1604 => to_slv(opcode_type, 16#0B#),
      1605 => to_slv(opcode_type, 16#08#),
      1606 => to_slv(opcode_type, 16#11#),
      1607 => to_slv(opcode_type, 16#0A#),
      1608 => to_slv(opcode_type, 16#06#),
      1609 => to_slv(opcode_type, 16#08#),
      1610 => to_slv(opcode_type, 16#03#),
      1611 => to_slv(opcode_type, 16#0A#),
      1612 => to_slv(opcode_type, 16#01#),
      1613 => to_slv(opcode_type, 16#0D#),
      1614 => to_slv(opcode_type, 16#07#),
      1615 => to_slv(opcode_type, 16#06#),
      1616 => to_slv(opcode_type, 16#0B#),
      1617 => to_slv(opcode_type, 16#32#),
      1618 => to_slv(opcode_type, 16#01#),
      1619 => to_slv(opcode_type, 16#0A#),
      1620 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#06#),
      1633 => to_slv(opcode_type, 16#07#),
      1634 => to_slv(opcode_type, 16#07#),
      1635 => to_slv(opcode_type, 16#06#),
      1636 => to_slv(opcode_type, 16#0D#),
      1637 => to_slv(opcode_type, 16#11#),
      1638 => to_slv(opcode_type, 16#05#),
      1639 => to_slv(opcode_type, 16#11#),
      1640 => to_slv(opcode_type, 16#06#),
      1641 => to_slv(opcode_type, 16#07#),
      1642 => to_slv(opcode_type, 16#0B#),
      1643 => to_slv(opcode_type, 16#0C#),
      1644 => to_slv(opcode_type, 16#07#),
      1645 => to_slv(opcode_type, 16#0C#),
      1646 => to_slv(opcode_type, 16#10#),
      1647 => to_slv(opcode_type, 16#05#),
      1648 => to_slv(opcode_type, 16#05#),
      1649 => to_slv(opcode_type, 16#07#),
      1650 => to_slv(opcode_type, 16#0E#),
      1651 => to_slv(opcode_type, 16#0F#),
      1652 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#08#),
      1665 => to_slv(opcode_type, 16#07#),
      1666 => to_slv(opcode_type, 16#07#),
      1667 => to_slv(opcode_type, 16#09#),
      1668 => to_slv(opcode_type, 16#0A#),
      1669 => to_slv(opcode_type, 16#0F#),
      1670 => to_slv(opcode_type, 16#05#),
      1671 => to_slv(opcode_type, 16#DB#),
      1672 => to_slv(opcode_type, 16#03#),
      1673 => to_slv(opcode_type, 16#02#),
      1674 => to_slv(opcode_type, 16#A6#),
      1675 => to_slv(opcode_type, 16#09#),
      1676 => to_slv(opcode_type, 16#07#),
      1677 => to_slv(opcode_type, 16#06#),
      1678 => to_slv(opcode_type, 16#0E#),
      1679 => to_slv(opcode_type, 16#10#),
      1680 => to_slv(opcode_type, 16#09#),
      1681 => to_slv(opcode_type, 16#0B#),
      1682 => to_slv(opcode_type, 16#68#),
      1683 => to_slv(opcode_type, 16#0C#),
      1684 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#06#),
      1697 => to_slv(opcode_type, 16#05#),
      1698 => to_slv(opcode_type, 16#08#),
      1699 => to_slv(opcode_type, 16#02#),
      1700 => to_slv(opcode_type, 16#0F#),
      1701 => to_slv(opcode_type, 16#05#),
      1702 => to_slv(opcode_type, 16#0F#),
      1703 => to_slv(opcode_type, 16#09#),
      1704 => to_slv(opcode_type, 16#08#),
      1705 => to_slv(opcode_type, 16#05#),
      1706 => to_slv(opcode_type, 16#0B#),
      1707 => to_slv(opcode_type, 16#09#),
      1708 => to_slv(opcode_type, 16#15#),
      1709 => to_slv(opcode_type, 16#0D#),
      1710 => to_slv(opcode_type, 16#07#),
      1711 => to_slv(opcode_type, 16#08#),
      1712 => to_slv(opcode_type, 16#0D#),
      1713 => to_slv(opcode_type, 16#0C#),
      1714 => to_slv(opcode_type, 16#02#),
      1715 => to_slv(opcode_type, 16#0A#),
      1716 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#08#),
      1729 => to_slv(opcode_type, 16#02#),
      1730 => to_slv(opcode_type, 16#02#),
      1731 => to_slv(opcode_type, 16#03#),
      1732 => to_slv(opcode_type, 16#11#),
      1733 => to_slv(opcode_type, 16#07#),
      1734 => to_slv(opcode_type, 16#07#),
      1735 => to_slv(opcode_type, 16#08#),
      1736 => to_slv(opcode_type, 16#0C#),
      1737 => to_slv(opcode_type, 16#11#),
      1738 => to_slv(opcode_type, 16#08#),
      1739 => to_slv(opcode_type, 16#0F#),
      1740 => to_slv(opcode_type, 16#0F#),
      1741 => to_slv(opcode_type, 16#09#),
      1742 => to_slv(opcode_type, 16#08#),
      1743 => to_slv(opcode_type, 16#0F#),
      1744 => to_slv(opcode_type, 16#0E#),
      1745 => to_slv(opcode_type, 16#07#),
      1746 => to_slv(opcode_type, 16#0F#),
      1747 => to_slv(opcode_type, 16#0D#),
      1748 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#06#),
      1761 => to_slv(opcode_type, 16#04#),
      1762 => to_slv(opcode_type, 16#09#),
      1763 => to_slv(opcode_type, 16#07#),
      1764 => to_slv(opcode_type, 16#10#),
      1765 => to_slv(opcode_type, 16#0B#),
      1766 => to_slv(opcode_type, 16#08#),
      1767 => to_slv(opcode_type, 16#0B#),
      1768 => to_slv(opcode_type, 16#0A#),
      1769 => to_slv(opcode_type, 16#07#),
      1770 => to_slv(opcode_type, 16#08#),
      1771 => to_slv(opcode_type, 16#08#),
      1772 => to_slv(opcode_type, 16#11#),
      1773 => to_slv(opcode_type, 16#0A#),
      1774 => to_slv(opcode_type, 16#08#),
      1775 => to_slv(opcode_type, 16#10#),
      1776 => to_slv(opcode_type, 16#11#),
      1777 => to_slv(opcode_type, 16#02#),
      1778 => to_slv(opcode_type, 16#04#),
      1779 => to_slv(opcode_type, 16#0A#),
      1780 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#06#),
      1793 => to_slv(opcode_type, 16#04#),
      1794 => to_slv(opcode_type, 16#09#),
      1795 => to_slv(opcode_type, 16#09#),
      1796 => to_slv(opcode_type, 16#0A#),
      1797 => to_slv(opcode_type, 16#10#),
      1798 => to_slv(opcode_type, 16#03#),
      1799 => to_slv(opcode_type, 16#0F#),
      1800 => to_slv(opcode_type, 16#09#),
      1801 => to_slv(opcode_type, 16#08#),
      1802 => to_slv(opcode_type, 16#01#),
      1803 => to_slv(opcode_type, 16#0B#),
      1804 => to_slv(opcode_type, 16#04#),
      1805 => to_slv(opcode_type, 16#0E#),
      1806 => to_slv(opcode_type, 16#08#),
      1807 => to_slv(opcode_type, 16#01#),
      1808 => to_slv(opcode_type, 16#0D#),
      1809 => to_slv(opcode_type, 16#06#),
      1810 => to_slv(opcode_type, 16#11#),
      1811 => to_slv(opcode_type, 16#0E#),
      1812 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#06#),
      1825 => to_slv(opcode_type, 16#04#),
      1826 => to_slv(opcode_type, 16#02#),
      1827 => to_slv(opcode_type, 16#04#),
      1828 => to_slv(opcode_type, 16#0A#),
      1829 => to_slv(opcode_type, 16#07#),
      1830 => to_slv(opcode_type, 16#09#),
      1831 => to_slv(opcode_type, 16#09#),
      1832 => to_slv(opcode_type, 16#0B#),
      1833 => to_slv(opcode_type, 16#0D#),
      1834 => to_slv(opcode_type, 16#08#),
      1835 => to_slv(opcode_type, 16#0F#),
      1836 => to_slv(opcode_type, 16#0C#),
      1837 => to_slv(opcode_type, 16#08#),
      1838 => to_slv(opcode_type, 16#06#),
      1839 => to_slv(opcode_type, 16#0B#),
      1840 => to_slv(opcode_type, 16#11#),
      1841 => to_slv(opcode_type, 16#08#),
      1842 => to_slv(opcode_type, 16#B7#),
      1843 => to_slv(opcode_type, 16#11#),
      1844 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#09#),
      1857 => to_slv(opcode_type, 16#04#),
      1858 => to_slv(opcode_type, 16#03#),
      1859 => to_slv(opcode_type, 16#08#),
      1860 => to_slv(opcode_type, 16#24#),
      1861 => to_slv(opcode_type, 16#F3#),
      1862 => to_slv(opcode_type, 16#07#),
      1863 => to_slv(opcode_type, 16#06#),
      1864 => to_slv(opcode_type, 16#05#),
      1865 => to_slv(opcode_type, 16#11#),
      1866 => to_slv(opcode_type, 16#07#),
      1867 => to_slv(opcode_type, 16#0E#),
      1868 => to_slv(opcode_type, 16#0C#),
      1869 => to_slv(opcode_type, 16#06#),
      1870 => to_slv(opcode_type, 16#07#),
      1871 => to_slv(opcode_type, 16#0B#),
      1872 => to_slv(opcode_type, 16#0E#),
      1873 => to_slv(opcode_type, 16#06#),
      1874 => to_slv(opcode_type, 16#0C#),
      1875 => to_slv(opcode_type, 16#0A#),
      1876 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#01#),
      1890 => to_slv(opcode_type, 16#01#),
      1891 => to_slv(opcode_type, 16#07#),
      1892 => to_slv(opcode_type, 16#0E#),
      1893 => to_slv(opcode_type, 16#10#),
      1894 => to_slv(opcode_type, 16#07#),
      1895 => to_slv(opcode_type, 16#07#),
      1896 => to_slv(opcode_type, 16#09#),
      1897 => to_slv(opcode_type, 16#0E#),
      1898 => to_slv(opcode_type, 16#0E#),
      1899 => to_slv(opcode_type, 16#03#),
      1900 => to_slv(opcode_type, 16#D7#),
      1901 => to_slv(opcode_type, 16#06#),
      1902 => to_slv(opcode_type, 16#06#),
      1903 => to_slv(opcode_type, 16#0C#),
      1904 => to_slv(opcode_type, 16#0B#),
      1905 => to_slv(opcode_type, 16#09#),
      1906 => to_slv(opcode_type, 16#0D#),
      1907 => to_slv(opcode_type, 16#0F#),
      1908 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#06#),
      1921 => to_slv(opcode_type, 16#07#),
      1922 => to_slv(opcode_type, 16#01#),
      1923 => to_slv(opcode_type, 16#01#),
      1924 => to_slv(opcode_type, 16#0F#),
      1925 => to_slv(opcode_type, 16#07#),
      1926 => to_slv(opcode_type, 16#08#),
      1927 => to_slv(opcode_type, 16#0A#),
      1928 => to_slv(opcode_type, 16#11#),
      1929 => to_slv(opcode_type, 16#08#),
      1930 => to_slv(opcode_type, 16#0C#),
      1931 => to_slv(opcode_type, 16#39#),
      1932 => to_slv(opcode_type, 16#08#),
      1933 => to_slv(opcode_type, 16#03#),
      1934 => to_slv(opcode_type, 16#05#),
      1935 => to_slv(opcode_type, 16#0F#),
      1936 => to_slv(opcode_type, 16#07#),
      1937 => to_slv(opcode_type, 16#03#),
      1938 => to_slv(opcode_type, 16#0C#),
      1939 => to_slv(opcode_type, 16#0E#),
      1940 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#08#),
      1953 => to_slv(opcode_type, 16#06#),
      1954 => to_slv(opcode_type, 16#03#),
      1955 => to_slv(opcode_type, 16#06#),
      1956 => to_slv(opcode_type, 16#9B#),
      1957 => to_slv(opcode_type, 16#0C#),
      1958 => to_slv(opcode_type, 16#07#),
      1959 => to_slv(opcode_type, 16#04#),
      1960 => to_slv(opcode_type, 16#11#),
      1961 => to_slv(opcode_type, 16#07#),
      1962 => to_slv(opcode_type, 16#0C#),
      1963 => to_slv(opcode_type, 16#0B#),
      1964 => to_slv(opcode_type, 16#09#),
      1965 => to_slv(opcode_type, 16#05#),
      1966 => to_slv(opcode_type, 16#06#),
      1967 => to_slv(opcode_type, 16#0A#),
      1968 => to_slv(opcode_type, 16#0A#),
      1969 => to_slv(opcode_type, 16#04#),
      1970 => to_slv(opcode_type, 16#04#),
      1971 => to_slv(opcode_type, 16#0D#),
      1972 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#08#),
      1985 => to_slv(opcode_type, 16#07#),
      1986 => to_slv(opcode_type, 16#03#),
      1987 => to_slv(opcode_type, 16#07#),
      1988 => to_slv(opcode_type, 16#0C#),
      1989 => to_slv(opcode_type, 16#0C#),
      1990 => to_slv(opcode_type, 16#04#),
      1991 => to_slv(opcode_type, 16#05#),
      1992 => to_slv(opcode_type, 16#0E#),
      1993 => to_slv(opcode_type, 16#08#),
      1994 => to_slv(opcode_type, 16#01#),
      1995 => to_slv(opcode_type, 16#03#),
      1996 => to_slv(opcode_type, 16#0F#),
      1997 => to_slv(opcode_type, 16#07#),
      1998 => to_slv(opcode_type, 16#08#),
      1999 => to_slv(opcode_type, 16#11#),
      2000 => to_slv(opcode_type, 16#CB#),
      2001 => to_slv(opcode_type, 16#07#),
      2002 => to_slv(opcode_type, 16#0F#),
      2003 => to_slv(opcode_type, 16#0D#),
      2004 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#07#),
      2017 => to_slv(opcode_type, 16#01#),
      2018 => to_slv(opcode_type, 16#04#),
      2019 => to_slv(opcode_type, 16#01#),
      2020 => to_slv(opcode_type, 16#0A#),
      2021 => to_slv(opcode_type, 16#07#),
      2022 => to_slv(opcode_type, 16#06#),
      2023 => to_slv(opcode_type, 16#06#),
      2024 => to_slv(opcode_type, 16#11#),
      2025 => to_slv(opcode_type, 16#0E#),
      2026 => to_slv(opcode_type, 16#09#),
      2027 => to_slv(opcode_type, 16#0E#),
      2028 => to_slv(opcode_type, 16#0D#),
      2029 => to_slv(opcode_type, 16#07#),
      2030 => to_slv(opcode_type, 16#06#),
      2031 => to_slv(opcode_type, 16#11#),
      2032 => to_slv(opcode_type, 16#0C#),
      2033 => to_slv(opcode_type, 16#09#),
      2034 => to_slv(opcode_type, 16#0F#),
      2035 => to_slv(opcode_type, 16#0C#),
      2036 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#06#),
      2049 => to_slv(opcode_type, 16#04#),
      2050 => to_slv(opcode_type, 16#01#),
      2051 => to_slv(opcode_type, 16#07#),
      2052 => to_slv(opcode_type, 16#0C#),
      2053 => to_slv(opcode_type, 16#0C#),
      2054 => to_slv(opcode_type, 16#09#),
      2055 => to_slv(opcode_type, 16#08#),
      2056 => to_slv(opcode_type, 16#03#),
      2057 => to_slv(opcode_type, 16#0B#),
      2058 => to_slv(opcode_type, 16#07#),
      2059 => to_slv(opcode_type, 16#0D#),
      2060 => to_slv(opcode_type, 16#11#),
      2061 => to_slv(opcode_type, 16#07#),
      2062 => to_slv(opcode_type, 16#08#),
      2063 => to_slv(opcode_type, 16#10#),
      2064 => to_slv(opcode_type, 16#0F#),
      2065 => to_slv(opcode_type, 16#08#),
      2066 => to_slv(opcode_type, 16#0A#),
      2067 => to_slv(opcode_type, 16#0C#),
      2068 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#07#),
      2081 => to_slv(opcode_type, 16#04#),
      2082 => to_slv(opcode_type, 16#04#),
      2083 => to_slv(opcode_type, 16#09#),
      2084 => to_slv(opcode_type, 16#0E#),
      2085 => to_slv(opcode_type, 16#0C#),
      2086 => to_slv(opcode_type, 16#07#),
      2087 => to_slv(opcode_type, 16#07#),
      2088 => to_slv(opcode_type, 16#08#),
      2089 => to_slv(opcode_type, 16#10#),
      2090 => to_slv(opcode_type, 16#0D#),
      2091 => to_slv(opcode_type, 16#05#),
      2092 => to_slv(opcode_type, 16#1C#),
      2093 => to_slv(opcode_type, 16#08#),
      2094 => to_slv(opcode_type, 16#06#),
      2095 => to_slv(opcode_type, 16#11#),
      2096 => to_slv(opcode_type, 16#10#),
      2097 => to_slv(opcode_type, 16#08#),
      2098 => to_slv(opcode_type, 16#0C#),
      2099 => to_slv(opcode_type, 16#0A#),
      2100 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#08#),
      2113 => to_slv(opcode_type, 16#06#),
      2114 => to_slv(opcode_type, 16#02#),
      2115 => to_slv(opcode_type, 16#02#),
      2116 => to_slv(opcode_type, 16#0B#),
      2117 => to_slv(opcode_type, 16#02#),
      2118 => to_slv(opcode_type, 16#06#),
      2119 => to_slv(opcode_type, 16#10#),
      2120 => to_slv(opcode_type, 16#10#),
      2121 => to_slv(opcode_type, 16#08#),
      2122 => to_slv(opcode_type, 16#06#),
      2123 => to_slv(opcode_type, 16#08#),
      2124 => to_slv(opcode_type, 16#0C#),
      2125 => to_slv(opcode_type, 16#0C#),
      2126 => to_slv(opcode_type, 16#03#),
      2127 => to_slv(opcode_type, 16#11#),
      2128 => to_slv(opcode_type, 16#03#),
      2129 => to_slv(opcode_type, 16#07#),
      2130 => to_slv(opcode_type, 16#0C#),
      2131 => to_slv(opcode_type, 16#0C#),
      2132 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#06#),
      2145 => to_slv(opcode_type, 16#02#),
      2146 => to_slv(opcode_type, 16#03#),
      2147 => to_slv(opcode_type, 16#02#),
      2148 => to_slv(opcode_type, 16#2E#),
      2149 => to_slv(opcode_type, 16#06#),
      2150 => to_slv(opcode_type, 16#08#),
      2151 => to_slv(opcode_type, 16#07#),
      2152 => to_slv(opcode_type, 16#11#),
      2153 => to_slv(opcode_type, 16#11#),
      2154 => to_slv(opcode_type, 16#08#),
      2155 => to_slv(opcode_type, 16#0B#),
      2156 => to_slv(opcode_type, 16#73#),
      2157 => to_slv(opcode_type, 16#09#),
      2158 => to_slv(opcode_type, 16#09#),
      2159 => to_slv(opcode_type, 16#0D#),
      2160 => to_slv(opcode_type, 16#0F#),
      2161 => to_slv(opcode_type, 16#07#),
      2162 => to_slv(opcode_type, 16#0D#),
      2163 => to_slv(opcode_type, 16#0E#),
      2164 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#08#),
      2177 => to_slv(opcode_type, 16#05#),
      2178 => to_slv(opcode_type, 16#09#),
      2179 => to_slv(opcode_type, 16#02#),
      2180 => to_slv(opcode_type, 16#10#),
      2181 => to_slv(opcode_type, 16#09#),
      2182 => to_slv(opcode_type, 16#0A#),
      2183 => to_slv(opcode_type, 16#0A#),
      2184 => to_slv(opcode_type, 16#07#),
      2185 => to_slv(opcode_type, 16#04#),
      2186 => to_slv(opcode_type, 16#07#),
      2187 => to_slv(opcode_type, 16#22#),
      2188 => to_slv(opcode_type, 16#11#),
      2189 => to_slv(opcode_type, 16#08#),
      2190 => to_slv(opcode_type, 16#08#),
      2191 => to_slv(opcode_type, 16#11#),
      2192 => to_slv(opcode_type, 16#10#),
      2193 => to_slv(opcode_type, 16#08#),
      2194 => to_slv(opcode_type, 16#11#),
      2195 => to_slv(opcode_type, 16#10#),
      2196 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#06#),
      2209 => to_slv(opcode_type, 16#02#),
      2210 => to_slv(opcode_type, 16#07#),
      2211 => to_slv(opcode_type, 16#09#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#0F#),
      2214 => to_slv(opcode_type, 16#05#),
      2215 => to_slv(opcode_type, 16#0D#),
      2216 => to_slv(opcode_type, 16#07#),
      2217 => to_slv(opcode_type, 16#06#),
      2218 => to_slv(opcode_type, 16#06#),
      2219 => to_slv(opcode_type, 16#CD#),
      2220 => to_slv(opcode_type, 16#0C#),
      2221 => to_slv(opcode_type, 16#07#),
      2222 => to_slv(opcode_type, 16#0B#),
      2223 => to_slv(opcode_type, 16#0D#),
      2224 => to_slv(opcode_type, 16#02#),
      2225 => to_slv(opcode_type, 16#06#),
      2226 => to_slv(opcode_type, 16#0B#),
      2227 => to_slv(opcode_type, 16#0C#),
      2228 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#09#),
      2241 => to_slv(opcode_type, 16#04#),
      2242 => to_slv(opcode_type, 16#07#),
      2243 => to_slv(opcode_type, 16#07#),
      2244 => to_slv(opcode_type, 16#11#),
      2245 => to_slv(opcode_type, 16#0B#),
      2246 => to_slv(opcode_type, 16#09#),
      2247 => to_slv(opcode_type, 16#10#),
      2248 => to_slv(opcode_type, 16#11#),
      2249 => to_slv(opcode_type, 16#09#),
      2250 => to_slv(opcode_type, 16#03#),
      2251 => to_slv(opcode_type, 16#05#),
      2252 => to_slv(opcode_type, 16#0F#),
      2253 => to_slv(opcode_type, 16#07#),
      2254 => to_slv(opcode_type, 16#06#),
      2255 => to_slv(opcode_type, 16#0F#),
      2256 => to_slv(opcode_type, 16#41#),
      2257 => to_slv(opcode_type, 16#07#),
      2258 => to_slv(opcode_type, 16#0D#),
      2259 => to_slv(opcode_type, 16#0C#),
      2260 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#06#),
      2273 => to_slv(opcode_type, 16#02#),
      2274 => to_slv(opcode_type, 16#09#),
      2275 => to_slv(opcode_type, 16#07#),
      2276 => to_slv(opcode_type, 16#0B#),
      2277 => to_slv(opcode_type, 16#0C#),
      2278 => to_slv(opcode_type, 16#06#),
      2279 => to_slv(opcode_type, 16#0E#),
      2280 => to_slv(opcode_type, 16#0F#),
      2281 => to_slv(opcode_type, 16#07#),
      2282 => to_slv(opcode_type, 16#03#),
      2283 => to_slv(opcode_type, 16#01#),
      2284 => to_slv(opcode_type, 16#0A#),
      2285 => to_slv(opcode_type, 16#06#),
      2286 => to_slv(opcode_type, 16#09#),
      2287 => to_slv(opcode_type, 16#0F#),
      2288 => to_slv(opcode_type, 16#11#),
      2289 => to_slv(opcode_type, 16#09#),
      2290 => to_slv(opcode_type, 16#10#),
      2291 => to_slv(opcode_type, 16#EB#),
      2292 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#06#),
      2305 => to_slv(opcode_type, 16#02#),
      2306 => to_slv(opcode_type, 16#07#),
      2307 => to_slv(opcode_type, 16#03#),
      2308 => to_slv(opcode_type, 16#11#),
      2309 => to_slv(opcode_type, 16#06#),
      2310 => to_slv(opcode_type, 16#0D#),
      2311 => to_slv(opcode_type, 16#10#),
      2312 => to_slv(opcode_type, 16#09#),
      2313 => to_slv(opcode_type, 16#03#),
      2314 => to_slv(opcode_type, 16#07#),
      2315 => to_slv(opcode_type, 16#0B#),
      2316 => to_slv(opcode_type, 16#10#),
      2317 => to_slv(opcode_type, 16#07#),
      2318 => to_slv(opcode_type, 16#09#),
      2319 => to_slv(opcode_type, 16#0B#),
      2320 => to_slv(opcode_type, 16#11#),
      2321 => to_slv(opcode_type, 16#08#),
      2322 => to_slv(opcode_type, 16#0F#),
      2323 => to_slv(opcode_type, 16#0D#),
      2324 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#07#),
      2337 => to_slv(opcode_type, 16#01#),
      2338 => to_slv(opcode_type, 16#07#),
      2339 => to_slv(opcode_type, 16#08#),
      2340 => to_slv(opcode_type, 16#11#),
      2341 => to_slv(opcode_type, 16#0B#),
      2342 => to_slv(opcode_type, 16#07#),
      2343 => to_slv(opcode_type, 16#0B#),
      2344 => to_slv(opcode_type, 16#10#),
      2345 => to_slv(opcode_type, 16#07#),
      2346 => to_slv(opcode_type, 16#09#),
      2347 => to_slv(opcode_type, 16#06#),
      2348 => to_slv(opcode_type, 16#11#),
      2349 => to_slv(opcode_type, 16#11#),
      2350 => to_slv(opcode_type, 16#04#),
      2351 => to_slv(opcode_type, 16#0E#),
      2352 => to_slv(opcode_type, 16#03#),
      2353 => to_slv(opcode_type, 16#09#),
      2354 => to_slv(opcode_type, 16#0C#),
      2355 => to_slv(opcode_type, 16#10#),
      2356 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#09#),
      2369 => to_slv(opcode_type, 16#08#),
      2370 => to_slv(opcode_type, 16#02#),
      2371 => to_slv(opcode_type, 16#05#),
      2372 => to_slv(opcode_type, 16#0B#),
      2373 => to_slv(opcode_type, 16#03#),
      2374 => to_slv(opcode_type, 16#05#),
      2375 => to_slv(opcode_type, 16#0D#),
      2376 => to_slv(opcode_type, 16#09#),
      2377 => to_slv(opcode_type, 16#09#),
      2378 => to_slv(opcode_type, 16#09#),
      2379 => to_slv(opcode_type, 16#0E#),
      2380 => to_slv(opcode_type, 16#11#),
      2381 => to_slv(opcode_type, 16#09#),
      2382 => to_slv(opcode_type, 16#10#),
      2383 => to_slv(opcode_type, 16#11#),
      2384 => to_slv(opcode_type, 16#01#),
      2385 => to_slv(opcode_type, 16#06#),
      2386 => to_slv(opcode_type, 16#13#),
      2387 => to_slv(opcode_type, 16#0C#),
      2388 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#08#),
      2401 => to_slv(opcode_type, 16#08#),
      2402 => to_slv(opcode_type, 16#06#),
      2403 => to_slv(opcode_type, 16#05#),
      2404 => to_slv(opcode_type, 16#11#),
      2405 => to_slv(opcode_type, 16#02#),
      2406 => to_slv(opcode_type, 16#0C#),
      2407 => to_slv(opcode_type, 16#06#),
      2408 => to_slv(opcode_type, 16#06#),
      2409 => to_slv(opcode_type, 16#0C#),
      2410 => to_slv(opcode_type, 16#A3#),
      2411 => to_slv(opcode_type, 16#06#),
      2412 => to_slv(opcode_type, 16#0B#),
      2413 => to_slv(opcode_type, 16#0A#),
      2414 => to_slv(opcode_type, 16#09#),
      2415 => to_slv(opcode_type, 16#05#),
      2416 => to_slv(opcode_type, 16#07#),
      2417 => to_slv(opcode_type, 16#7E#),
      2418 => to_slv(opcode_type, 16#10#),
      2419 => to_slv(opcode_type, 16#0E#),
      2420 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#08#),
      2433 => to_slv(opcode_type, 16#09#),
      2434 => to_slv(opcode_type, 16#04#),
      2435 => to_slv(opcode_type, 16#08#),
      2436 => to_slv(opcode_type, 16#3C#),
      2437 => to_slv(opcode_type, 16#10#),
      2438 => to_slv(opcode_type, 16#07#),
      2439 => to_slv(opcode_type, 16#09#),
      2440 => to_slv(opcode_type, 16#10#),
      2441 => to_slv(opcode_type, 16#0F#),
      2442 => to_slv(opcode_type, 16#09#),
      2443 => to_slv(opcode_type, 16#0D#),
      2444 => to_slv(opcode_type, 16#0C#),
      2445 => to_slv(opcode_type, 16#01#),
      2446 => to_slv(opcode_type, 16#09#),
      2447 => to_slv(opcode_type, 16#05#),
      2448 => to_slv(opcode_type, 16#0B#),
      2449 => to_slv(opcode_type, 16#09#),
      2450 => to_slv(opcode_type, 16#0F#),
      2451 => to_slv(opcode_type, 16#0A#),
      2452 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#09#),
      2465 => to_slv(opcode_type, 16#03#),
      2466 => to_slv(opcode_type, 16#08#),
      2467 => to_slv(opcode_type, 16#03#),
      2468 => to_slv(opcode_type, 16#0A#),
      2469 => to_slv(opcode_type, 16#07#),
      2470 => to_slv(opcode_type, 16#0A#),
      2471 => to_slv(opcode_type, 16#0E#),
      2472 => to_slv(opcode_type, 16#08#),
      2473 => to_slv(opcode_type, 16#03#),
      2474 => to_slv(opcode_type, 16#08#),
      2475 => to_slv(opcode_type, 16#4D#),
      2476 => to_slv(opcode_type, 16#10#),
      2477 => to_slv(opcode_type, 16#09#),
      2478 => to_slv(opcode_type, 16#06#),
      2479 => to_slv(opcode_type, 16#11#),
      2480 => to_slv(opcode_type, 16#0C#),
      2481 => to_slv(opcode_type, 16#06#),
      2482 => to_slv(opcode_type, 16#0D#),
      2483 => to_slv(opcode_type, 16#0C#),
      2484 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#07#),
      2497 => to_slv(opcode_type, 16#02#),
      2498 => to_slv(opcode_type, 16#03#),
      2499 => to_slv(opcode_type, 16#07#),
      2500 => to_slv(opcode_type, 16#0C#),
      2501 => to_slv(opcode_type, 16#10#),
      2502 => to_slv(opcode_type, 16#09#),
      2503 => to_slv(opcode_type, 16#07#),
      2504 => to_slv(opcode_type, 16#08#),
      2505 => to_slv(opcode_type, 16#0E#),
      2506 => to_slv(opcode_type, 16#0E#),
      2507 => to_slv(opcode_type, 16#01#),
      2508 => to_slv(opcode_type, 16#0F#),
      2509 => to_slv(opcode_type, 16#07#),
      2510 => to_slv(opcode_type, 16#09#),
      2511 => to_slv(opcode_type, 16#0C#),
      2512 => to_slv(opcode_type, 16#10#),
      2513 => to_slv(opcode_type, 16#09#),
      2514 => to_slv(opcode_type, 16#10#),
      2515 => to_slv(opcode_type, 16#10#),
      2516 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#07#),
      2530 => to_slv(opcode_type, 16#06#),
      2531 => to_slv(opcode_type, 16#06#),
      2532 => to_slv(opcode_type, 16#0D#),
      2533 => to_slv(opcode_type, 16#0A#),
      2534 => to_slv(opcode_type, 16#03#),
      2535 => to_slv(opcode_type, 16#82#),
      2536 => to_slv(opcode_type, 16#08#),
      2537 => to_slv(opcode_type, 16#01#),
      2538 => to_slv(opcode_type, 16#0B#),
      2539 => to_slv(opcode_type, 16#03#),
      2540 => to_slv(opcode_type, 16#0F#),
      2541 => to_slv(opcode_type, 16#05#),
      2542 => to_slv(opcode_type, 16#07#),
      2543 => to_slv(opcode_type, 16#07#),
      2544 => to_slv(opcode_type, 16#0F#),
      2545 => to_slv(opcode_type, 16#0F#),
      2546 => to_slv(opcode_type, 16#03#),
      2547 => to_slv(opcode_type, 16#0F#),
      2548 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#09#),
      2561 => to_slv(opcode_type, 16#01#),
      2562 => to_slv(opcode_type, 16#03#),
      2563 => to_slv(opcode_type, 16#02#),
      2564 => to_slv(opcode_type, 16#0F#),
      2565 => to_slv(opcode_type, 16#09#),
      2566 => to_slv(opcode_type, 16#06#),
      2567 => to_slv(opcode_type, 16#06#),
      2568 => to_slv(opcode_type, 16#0A#),
      2569 => to_slv(opcode_type, 16#0F#),
      2570 => to_slv(opcode_type, 16#08#),
      2571 => to_slv(opcode_type, 16#0F#),
      2572 => to_slv(opcode_type, 16#0A#),
      2573 => to_slv(opcode_type, 16#09#),
      2574 => to_slv(opcode_type, 16#08#),
      2575 => to_slv(opcode_type, 16#0B#),
      2576 => to_slv(opcode_type, 16#0E#),
      2577 => to_slv(opcode_type, 16#08#),
      2578 => to_slv(opcode_type, 16#10#),
      2579 => to_slv(opcode_type, 16#0F#),
      2580 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#08#),
      2593 => to_slv(opcode_type, 16#09#),
      2594 => to_slv(opcode_type, 16#03#),
      2595 => to_slv(opcode_type, 16#08#),
      2596 => to_slv(opcode_type, 16#0C#),
      2597 => to_slv(opcode_type, 16#0B#),
      2598 => to_slv(opcode_type, 16#04#),
      2599 => to_slv(opcode_type, 16#02#),
      2600 => to_slv(opcode_type, 16#0A#),
      2601 => to_slv(opcode_type, 16#09#),
      2602 => to_slv(opcode_type, 16#03#),
      2603 => to_slv(opcode_type, 16#09#),
      2604 => to_slv(opcode_type, 16#10#),
      2605 => to_slv(opcode_type, 16#E3#),
      2606 => to_slv(opcode_type, 16#06#),
      2607 => to_slv(opcode_type, 16#05#),
      2608 => to_slv(opcode_type, 16#0C#),
      2609 => to_slv(opcode_type, 16#06#),
      2610 => to_slv(opcode_type, 16#10#),
      2611 => to_slv(opcode_type, 16#0A#),
      2612 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#09#),
      2625 => to_slv(opcode_type, 16#05#),
      2626 => to_slv(opcode_type, 16#07#),
      2627 => to_slv(opcode_type, 16#06#),
      2628 => to_slv(opcode_type, 16#0C#),
      2629 => to_slv(opcode_type, 16#0F#),
      2630 => to_slv(opcode_type, 16#05#),
      2631 => to_slv(opcode_type, 16#0E#),
      2632 => to_slv(opcode_type, 16#08#),
      2633 => to_slv(opcode_type, 16#05#),
      2634 => to_slv(opcode_type, 16#07#),
      2635 => to_slv(opcode_type, 16#0F#),
      2636 => to_slv(opcode_type, 16#10#),
      2637 => to_slv(opcode_type, 16#07#),
      2638 => to_slv(opcode_type, 16#08#),
      2639 => to_slv(opcode_type, 16#0C#),
      2640 => to_slv(opcode_type, 16#DB#),
      2641 => to_slv(opcode_type, 16#09#),
      2642 => to_slv(opcode_type, 16#0A#),
      2643 => to_slv(opcode_type, 16#10#),
      2644 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#07#),
      2657 => to_slv(opcode_type, 16#07#),
      2658 => to_slv(opcode_type, 16#09#),
      2659 => to_slv(opcode_type, 16#07#),
      2660 => to_slv(opcode_type, 16#0E#),
      2661 => to_slv(opcode_type, 16#0D#),
      2662 => to_slv(opcode_type, 16#06#),
      2663 => to_slv(opcode_type, 16#10#),
      2664 => to_slv(opcode_type, 16#0F#),
      2665 => to_slv(opcode_type, 16#03#),
      2666 => to_slv(opcode_type, 16#06#),
      2667 => to_slv(opcode_type, 16#0F#),
      2668 => to_slv(opcode_type, 16#10#),
      2669 => to_slv(opcode_type, 16#02#),
      2670 => to_slv(opcode_type, 16#07#),
      2671 => to_slv(opcode_type, 16#08#),
      2672 => to_slv(opcode_type, 16#0A#),
      2673 => to_slv(opcode_type, 16#10#),
      2674 => to_slv(opcode_type, 16#01#),
      2675 => to_slv(opcode_type, 16#0F#),
      2676 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#09#),
      2689 => to_slv(opcode_type, 16#05#),
      2690 => to_slv(opcode_type, 16#04#),
      2691 => to_slv(opcode_type, 16#05#),
      2692 => to_slv(opcode_type, 16#0C#),
      2693 => to_slv(opcode_type, 16#06#),
      2694 => to_slv(opcode_type, 16#09#),
      2695 => to_slv(opcode_type, 16#07#),
      2696 => to_slv(opcode_type, 16#0E#),
      2697 => to_slv(opcode_type, 16#0E#),
      2698 => to_slv(opcode_type, 16#06#),
      2699 => to_slv(opcode_type, 16#0C#),
      2700 => to_slv(opcode_type, 16#0F#),
      2701 => to_slv(opcode_type, 16#08#),
      2702 => to_slv(opcode_type, 16#06#),
      2703 => to_slv(opcode_type, 16#0A#),
      2704 => to_slv(opcode_type, 16#0A#),
      2705 => to_slv(opcode_type, 16#08#),
      2706 => to_slv(opcode_type, 16#0E#),
      2707 => to_slv(opcode_type, 16#0C#),
      2708 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#08#),
      2721 => to_slv(opcode_type, 16#08#),
      2722 => to_slv(opcode_type, 16#03#),
      2723 => to_slv(opcode_type, 16#04#),
      2724 => to_slv(opcode_type, 16#0B#),
      2725 => to_slv(opcode_type, 16#07#),
      2726 => to_slv(opcode_type, 16#03#),
      2727 => to_slv(opcode_type, 16#11#),
      2728 => to_slv(opcode_type, 16#08#),
      2729 => to_slv(opcode_type, 16#10#),
      2730 => to_slv(opcode_type, 16#0B#),
      2731 => to_slv(opcode_type, 16#07#),
      2732 => to_slv(opcode_type, 16#07#),
      2733 => to_slv(opcode_type, 16#07#),
      2734 => to_slv(opcode_type, 16#0A#),
      2735 => to_slv(opcode_type, 16#0E#),
      2736 => to_slv(opcode_type, 16#03#),
      2737 => to_slv(opcode_type, 16#10#),
      2738 => to_slv(opcode_type, 16#04#),
      2739 => to_slv(opcode_type, 16#10#),
      2740 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#07#),
      2753 => to_slv(opcode_type, 16#05#),
      2754 => to_slv(opcode_type, 16#06#),
      2755 => to_slv(opcode_type, 16#08#),
      2756 => to_slv(opcode_type, 16#0D#),
      2757 => to_slv(opcode_type, 16#0C#),
      2758 => to_slv(opcode_type, 16#03#),
      2759 => to_slv(opcode_type, 16#0A#),
      2760 => to_slv(opcode_type, 16#07#),
      2761 => to_slv(opcode_type, 16#08#),
      2762 => to_slv(opcode_type, 16#07#),
      2763 => to_slv(opcode_type, 16#CD#),
      2764 => to_slv(opcode_type, 16#0C#),
      2765 => to_slv(opcode_type, 16#04#),
      2766 => to_slv(opcode_type, 16#0C#),
      2767 => to_slv(opcode_type, 16#09#),
      2768 => to_slv(opcode_type, 16#05#),
      2769 => to_slv(opcode_type, 16#DF#),
      2770 => to_slv(opcode_type, 16#01#),
      2771 => to_slv(opcode_type, 16#0F#),
      2772 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#07#),
      2785 => to_slv(opcode_type, 16#03#),
      2786 => to_slv(opcode_type, 16#03#),
      2787 => to_slv(opcode_type, 16#01#),
      2788 => to_slv(opcode_type, 16#0C#),
      2789 => to_slv(opcode_type, 16#07#),
      2790 => to_slv(opcode_type, 16#07#),
      2791 => to_slv(opcode_type, 16#07#),
      2792 => to_slv(opcode_type, 16#0C#),
      2793 => to_slv(opcode_type, 16#0C#),
      2794 => to_slv(opcode_type, 16#08#),
      2795 => to_slv(opcode_type, 16#11#),
      2796 => to_slv(opcode_type, 16#0B#),
      2797 => to_slv(opcode_type, 16#09#),
      2798 => to_slv(opcode_type, 16#08#),
      2799 => to_slv(opcode_type, 16#0C#),
      2800 => to_slv(opcode_type, 16#11#),
      2801 => to_slv(opcode_type, 16#09#),
      2802 => to_slv(opcode_type, 16#10#),
      2803 => to_slv(opcode_type, 16#0E#),
      2804 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#08#),
      2817 => to_slv(opcode_type, 16#04#),
      2818 => to_slv(opcode_type, 16#07#),
      2819 => to_slv(opcode_type, 16#04#),
      2820 => to_slv(opcode_type, 16#0E#),
      2821 => to_slv(opcode_type, 16#01#),
      2822 => to_slv(opcode_type, 16#0F#),
      2823 => to_slv(opcode_type, 16#08#),
      2824 => to_slv(opcode_type, 16#07#),
      2825 => to_slv(opcode_type, 16#03#),
      2826 => to_slv(opcode_type, 16#0B#),
      2827 => to_slv(opcode_type, 16#08#),
      2828 => to_slv(opcode_type, 16#0C#),
      2829 => to_slv(opcode_type, 16#10#),
      2830 => to_slv(opcode_type, 16#09#),
      2831 => to_slv(opcode_type, 16#04#),
      2832 => to_slv(opcode_type, 16#0F#),
      2833 => to_slv(opcode_type, 16#08#),
      2834 => to_slv(opcode_type, 16#10#),
      2835 => to_slv(opcode_type, 16#11#),
      2836 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#08#),
      2849 => to_slv(opcode_type, 16#09#),
      2850 => to_slv(opcode_type, 16#08#),
      2851 => to_slv(opcode_type, 16#07#),
      2852 => to_slv(opcode_type, 16#10#),
      2853 => to_slv(opcode_type, 16#11#),
      2854 => to_slv(opcode_type, 16#04#),
      2855 => to_slv(opcode_type, 16#0D#),
      2856 => to_slv(opcode_type, 16#04#),
      2857 => to_slv(opcode_type, 16#04#),
      2858 => to_slv(opcode_type, 16#0B#),
      2859 => to_slv(opcode_type, 16#06#),
      2860 => to_slv(opcode_type, 16#08#),
      2861 => to_slv(opcode_type, 16#02#),
      2862 => to_slv(opcode_type, 16#0B#),
      2863 => to_slv(opcode_type, 16#08#),
      2864 => to_slv(opcode_type, 16#0B#),
      2865 => to_slv(opcode_type, 16#0E#),
      2866 => to_slv(opcode_type, 16#04#),
      2867 => to_slv(opcode_type, 16#0E#),
      2868 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#06#),
      2881 => to_slv(opcode_type, 16#05#),
      2882 => to_slv(opcode_type, 16#01#),
      2883 => to_slv(opcode_type, 16#01#),
      2884 => to_slv(opcode_type, 16#0C#),
      2885 => to_slv(opcode_type, 16#06#),
      2886 => to_slv(opcode_type, 16#08#),
      2887 => to_slv(opcode_type, 16#07#),
      2888 => to_slv(opcode_type, 16#0F#),
      2889 => to_slv(opcode_type, 16#0D#),
      2890 => to_slv(opcode_type, 16#08#),
      2891 => to_slv(opcode_type, 16#0D#),
      2892 => to_slv(opcode_type, 16#7C#),
      2893 => to_slv(opcode_type, 16#06#),
      2894 => to_slv(opcode_type, 16#09#),
      2895 => to_slv(opcode_type, 16#0E#),
      2896 => to_slv(opcode_type, 16#DE#),
      2897 => to_slv(opcode_type, 16#08#),
      2898 => to_slv(opcode_type, 16#10#),
      2899 => to_slv(opcode_type, 16#11#),
      2900 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#08#),
      2913 => to_slv(opcode_type, 16#01#),
      2914 => to_slv(opcode_type, 16#09#),
      2915 => to_slv(opcode_type, 16#09#),
      2916 => to_slv(opcode_type, 16#0E#),
      2917 => to_slv(opcode_type, 16#0C#),
      2918 => to_slv(opcode_type, 16#05#),
      2919 => to_slv(opcode_type, 16#0B#),
      2920 => to_slv(opcode_type, 16#06#),
      2921 => to_slv(opcode_type, 16#09#),
      2922 => to_slv(opcode_type, 16#01#),
      2923 => to_slv(opcode_type, 16#0B#),
      2924 => to_slv(opcode_type, 16#08#),
      2925 => to_slv(opcode_type, 16#10#),
      2926 => to_slv(opcode_type, 16#0E#),
      2927 => to_slv(opcode_type, 16#08#),
      2928 => to_slv(opcode_type, 16#09#),
      2929 => to_slv(opcode_type, 16#10#),
      2930 => to_slv(opcode_type, 16#0F#),
      2931 => to_slv(opcode_type, 16#0E#),
      2932 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#07#),
      2945 => to_slv(opcode_type, 16#07#),
      2946 => to_slv(opcode_type, 16#03#),
      2947 => to_slv(opcode_type, 16#01#),
      2948 => to_slv(opcode_type, 16#0A#),
      2949 => to_slv(opcode_type, 16#01#),
      2950 => to_slv(opcode_type, 16#06#),
      2951 => to_slv(opcode_type, 16#0D#),
      2952 => to_slv(opcode_type, 16#10#),
      2953 => to_slv(opcode_type, 16#08#),
      2954 => to_slv(opcode_type, 16#08#),
      2955 => to_slv(opcode_type, 16#03#),
      2956 => to_slv(opcode_type, 16#10#),
      2957 => to_slv(opcode_type, 16#06#),
      2958 => to_slv(opcode_type, 16#0D#),
      2959 => to_slv(opcode_type, 16#10#),
      2960 => to_slv(opcode_type, 16#06#),
      2961 => to_slv(opcode_type, 16#01#),
      2962 => to_slv(opcode_type, 16#0D#),
      2963 => to_slv(opcode_type, 16#0A#),
      2964 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#07#),
      2977 => to_slv(opcode_type, 16#06#),
      2978 => to_slv(opcode_type, 16#09#),
      2979 => to_slv(opcode_type, 16#06#),
      2980 => to_slv(opcode_type, 16#0E#),
      2981 => to_slv(opcode_type, 16#11#),
      2982 => to_slv(opcode_type, 16#07#),
      2983 => to_slv(opcode_type, 16#9F#),
      2984 => to_slv(opcode_type, 16#10#),
      2985 => to_slv(opcode_type, 16#04#),
      2986 => to_slv(opcode_type, 16#09#),
      2987 => to_slv(opcode_type, 16#0B#),
      2988 => to_slv(opcode_type, 16#FF#),
      2989 => to_slv(opcode_type, 16#06#),
      2990 => to_slv(opcode_type, 16#03#),
      2991 => to_slv(opcode_type, 16#02#),
      2992 => to_slv(opcode_type, 16#0F#),
      2993 => to_slv(opcode_type, 16#01#),
      2994 => to_slv(opcode_type, 16#01#),
      2995 => to_slv(opcode_type, 16#0A#),
      2996 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#06#),
      3009 => to_slv(opcode_type, 16#04#),
      3010 => to_slv(opcode_type, 16#06#),
      3011 => to_slv(opcode_type, 16#08#),
      3012 => to_slv(opcode_type, 16#0F#),
      3013 => to_slv(opcode_type, 16#0F#),
      3014 => to_slv(opcode_type, 16#08#),
      3015 => to_slv(opcode_type, 16#91#),
      3016 => to_slv(opcode_type, 16#10#),
      3017 => to_slv(opcode_type, 16#08#),
      3018 => to_slv(opcode_type, 16#08#),
      3019 => to_slv(opcode_type, 16#03#),
      3020 => to_slv(opcode_type, 16#0C#),
      3021 => to_slv(opcode_type, 16#03#),
      3022 => to_slv(opcode_type, 16#0C#),
      3023 => to_slv(opcode_type, 16#06#),
      3024 => to_slv(opcode_type, 16#05#),
      3025 => to_slv(opcode_type, 16#10#),
      3026 => to_slv(opcode_type, 16#03#),
      3027 => to_slv(opcode_type, 16#0C#),
      3028 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#06#),
      3041 => to_slv(opcode_type, 16#02#),
      3042 => to_slv(opcode_type, 16#06#),
      3043 => to_slv(opcode_type, 16#05#),
      3044 => to_slv(opcode_type, 16#0B#),
      3045 => to_slv(opcode_type, 16#08#),
      3046 => to_slv(opcode_type, 16#0B#),
      3047 => to_slv(opcode_type, 16#0C#),
      3048 => to_slv(opcode_type, 16#09#),
      3049 => to_slv(opcode_type, 16#08#),
      3050 => to_slv(opcode_type, 16#07#),
      3051 => to_slv(opcode_type, 16#0E#),
      3052 => to_slv(opcode_type, 16#0A#),
      3053 => to_slv(opcode_type, 16#01#),
      3054 => to_slv(opcode_type, 16#10#),
      3055 => to_slv(opcode_type, 16#08#),
      3056 => to_slv(opcode_type, 16#01#),
      3057 => to_slv(opcode_type, 16#0C#),
      3058 => to_slv(opcode_type, 16#02#),
      3059 => to_slv(opcode_type, 16#10#),
      3060 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#07#),
      3073 => to_slv(opcode_type, 16#04#),
      3074 => to_slv(opcode_type, 16#06#),
      3075 => to_slv(opcode_type, 16#08#),
      3076 => to_slv(opcode_type, 16#BF#),
      3077 => to_slv(opcode_type, 16#0C#),
      3078 => to_slv(opcode_type, 16#06#),
      3079 => to_slv(opcode_type, 16#10#),
      3080 => to_slv(opcode_type, 16#11#),
      3081 => to_slv(opcode_type, 16#06#),
      3082 => to_slv(opcode_type, 16#03#),
      3083 => to_slv(opcode_type, 16#09#),
      3084 => to_slv(opcode_type, 16#0C#),
      3085 => to_slv(opcode_type, 16#0D#),
      3086 => to_slv(opcode_type, 16#09#),
      3087 => to_slv(opcode_type, 16#05#),
      3088 => to_slv(opcode_type, 16#0E#),
      3089 => to_slv(opcode_type, 16#08#),
      3090 => to_slv(opcode_type, 16#0F#),
      3091 => to_slv(opcode_type, 16#0C#),
      3092 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#09#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#09#),
      3107 => to_slv(opcode_type, 16#01#),
      3108 => to_slv(opcode_type, 16#0B#),
      3109 => to_slv(opcode_type, 16#02#),
      3110 => to_slv(opcode_type, 16#0E#),
      3111 => to_slv(opcode_type, 16#05#),
      3112 => to_slv(opcode_type, 16#05#),
      3113 => to_slv(opcode_type, 16#0E#),
      3114 => to_slv(opcode_type, 16#07#),
      3115 => to_slv(opcode_type, 16#06#),
      3116 => to_slv(opcode_type, 16#07#),
      3117 => to_slv(opcode_type, 16#10#),
      3118 => to_slv(opcode_type, 16#0D#),
      3119 => to_slv(opcode_type, 16#08#),
      3120 => to_slv(opcode_type, 16#0B#),
      3121 => to_slv(opcode_type, 16#0C#),
      3122 => to_slv(opcode_type, 16#02#),
      3123 => to_slv(opcode_type, 16#0F#),
      3124 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#06#),
      3137 => to_slv(opcode_type, 16#05#),
      3138 => to_slv(opcode_type, 16#06#),
      3139 => to_slv(opcode_type, 16#05#),
      3140 => to_slv(opcode_type, 16#0A#),
      3141 => to_slv(opcode_type, 16#02#),
      3142 => to_slv(opcode_type, 16#0F#),
      3143 => to_slv(opcode_type, 16#06#),
      3144 => to_slv(opcode_type, 16#08#),
      3145 => to_slv(opcode_type, 16#08#),
      3146 => to_slv(opcode_type, 16#0D#),
      3147 => to_slv(opcode_type, 16#11#),
      3148 => to_slv(opcode_type, 16#01#),
      3149 => to_slv(opcode_type, 16#0F#),
      3150 => to_slv(opcode_type, 16#09#),
      3151 => to_slv(opcode_type, 16#09#),
      3152 => to_slv(opcode_type, 16#0C#),
      3153 => to_slv(opcode_type, 16#0E#),
      3154 => to_slv(opcode_type, 16#03#),
      3155 => to_slv(opcode_type, 16#0B#),
      3156 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#06#),
      3169 => to_slv(opcode_type, 16#07#),
      3170 => to_slv(opcode_type, 16#01#),
      3171 => to_slv(opcode_type, 16#06#),
      3172 => to_slv(opcode_type, 16#0B#),
      3173 => to_slv(opcode_type, 16#0D#),
      3174 => to_slv(opcode_type, 16#05#),
      3175 => to_slv(opcode_type, 16#09#),
      3176 => to_slv(opcode_type, 16#16#),
      3177 => to_slv(opcode_type, 16#2B#),
      3178 => to_slv(opcode_type, 16#06#),
      3179 => to_slv(opcode_type, 16#03#),
      3180 => to_slv(opcode_type, 16#03#),
      3181 => to_slv(opcode_type, 16#0A#),
      3182 => to_slv(opcode_type, 16#09#),
      3183 => to_slv(opcode_type, 16#04#),
      3184 => to_slv(opcode_type, 16#0F#),
      3185 => to_slv(opcode_type, 16#07#),
      3186 => to_slv(opcode_type, 16#4D#),
      3187 => to_slv(opcode_type, 16#0D#),
      3188 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#07#),
      3201 => to_slv(opcode_type, 16#08#),
      3202 => to_slv(opcode_type, 16#01#),
      3203 => to_slv(opcode_type, 16#08#),
      3204 => to_slv(opcode_type, 16#0F#),
      3205 => to_slv(opcode_type, 16#0F#),
      3206 => to_slv(opcode_type, 16#06#),
      3207 => to_slv(opcode_type, 16#06#),
      3208 => to_slv(opcode_type, 16#0D#),
      3209 => to_slv(opcode_type, 16#0D#),
      3210 => to_slv(opcode_type, 16#02#),
      3211 => to_slv(opcode_type, 16#0B#),
      3212 => to_slv(opcode_type, 16#07#),
      3213 => to_slv(opcode_type, 16#09#),
      3214 => to_slv(opcode_type, 16#06#),
      3215 => to_slv(opcode_type, 16#0B#),
      3216 => to_slv(opcode_type, 16#0C#),
      3217 => to_slv(opcode_type, 16#02#),
      3218 => to_slv(opcode_type, 16#0F#),
      3219 => to_slv(opcode_type, 16#0B#),
      3220 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#09#),
      3233 => to_slv(opcode_type, 16#03#),
      3234 => to_slv(opcode_type, 16#01#),
      3235 => to_slv(opcode_type, 16#01#),
      3236 => to_slv(opcode_type, 16#11#),
      3237 => to_slv(opcode_type, 16#06#),
      3238 => to_slv(opcode_type, 16#09#),
      3239 => to_slv(opcode_type, 16#06#),
      3240 => to_slv(opcode_type, 16#0E#),
      3241 => to_slv(opcode_type, 16#C0#),
      3242 => to_slv(opcode_type, 16#07#),
      3243 => to_slv(opcode_type, 16#0A#),
      3244 => to_slv(opcode_type, 16#0C#),
      3245 => to_slv(opcode_type, 16#06#),
      3246 => to_slv(opcode_type, 16#09#),
      3247 => to_slv(opcode_type, 16#66#),
      3248 => to_slv(opcode_type, 16#0F#),
      3249 => to_slv(opcode_type, 16#06#),
      3250 => to_slv(opcode_type, 16#0C#),
      3251 => to_slv(opcode_type, 16#10#),
      3252 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#07#),
      3265 => to_slv(opcode_type, 16#07#),
      3266 => to_slv(opcode_type, 16#03#),
      3267 => to_slv(opcode_type, 16#04#),
      3268 => to_slv(opcode_type, 16#0C#),
      3269 => to_slv(opcode_type, 16#07#),
      3270 => to_slv(opcode_type, 16#07#),
      3271 => to_slv(opcode_type, 16#A1#),
      3272 => to_slv(opcode_type, 16#11#),
      3273 => to_slv(opcode_type, 16#08#),
      3274 => to_slv(opcode_type, 16#0C#),
      3275 => to_slv(opcode_type, 16#0D#),
      3276 => to_slv(opcode_type, 16#09#),
      3277 => to_slv(opcode_type, 16#04#),
      3278 => to_slv(opcode_type, 16#04#),
      3279 => to_slv(opcode_type, 16#B1#),
      3280 => to_slv(opcode_type, 16#06#),
      3281 => to_slv(opcode_type, 16#05#),
      3282 => to_slv(opcode_type, 16#11#),
      3283 => to_slv(opcode_type, 16#0A#),
      3284 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#06#),
      3297 => to_slv(opcode_type, 16#01#),
      3298 => to_slv(opcode_type, 16#03#),
      3299 => to_slv(opcode_type, 16#08#),
      3300 => to_slv(opcode_type, 16#0E#),
      3301 => to_slv(opcode_type, 16#D0#),
      3302 => to_slv(opcode_type, 16#06#),
      3303 => to_slv(opcode_type, 16#09#),
      3304 => to_slv(opcode_type, 16#04#),
      3305 => to_slv(opcode_type, 16#11#),
      3306 => to_slv(opcode_type, 16#08#),
      3307 => to_slv(opcode_type, 16#0A#),
      3308 => to_slv(opcode_type, 16#11#),
      3309 => to_slv(opcode_type, 16#08#),
      3310 => to_slv(opcode_type, 16#06#),
      3311 => to_slv(opcode_type, 16#10#),
      3312 => to_slv(opcode_type, 16#0A#),
      3313 => to_slv(opcode_type, 16#09#),
      3314 => to_slv(opcode_type, 16#11#),
      3315 => to_slv(opcode_type, 16#11#),
      3316 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#06#),
      3329 => to_slv(opcode_type, 16#08#),
      3330 => to_slv(opcode_type, 16#01#),
      3331 => to_slv(opcode_type, 16#08#),
      3332 => to_slv(opcode_type, 16#0D#),
      3333 => to_slv(opcode_type, 16#0E#),
      3334 => to_slv(opcode_type, 16#01#),
      3335 => to_slv(opcode_type, 16#05#),
      3336 => to_slv(opcode_type, 16#0B#),
      3337 => to_slv(opcode_type, 16#07#),
      3338 => to_slv(opcode_type, 16#05#),
      3339 => to_slv(opcode_type, 16#04#),
      3340 => to_slv(opcode_type, 16#10#),
      3341 => to_slv(opcode_type, 16#08#),
      3342 => to_slv(opcode_type, 16#06#),
      3343 => to_slv(opcode_type, 16#0B#),
      3344 => to_slv(opcode_type, 16#0B#),
      3345 => to_slv(opcode_type, 16#08#),
      3346 => to_slv(opcode_type, 16#F4#),
      3347 => to_slv(opcode_type, 16#11#),
      3348 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#09#),
      3361 => to_slv(opcode_type, 16#05#),
      3362 => to_slv(opcode_type, 16#03#),
      3363 => to_slv(opcode_type, 16#01#),
      3364 => to_slv(opcode_type, 16#0F#),
      3365 => to_slv(opcode_type, 16#09#),
      3366 => to_slv(opcode_type, 16#09#),
      3367 => to_slv(opcode_type, 16#06#),
      3368 => to_slv(opcode_type, 16#0A#),
      3369 => to_slv(opcode_type, 16#10#),
      3370 => to_slv(opcode_type, 16#07#),
      3371 => to_slv(opcode_type, 16#10#),
      3372 => to_slv(opcode_type, 16#0E#),
      3373 => to_slv(opcode_type, 16#08#),
      3374 => to_slv(opcode_type, 16#08#),
      3375 => to_slv(opcode_type, 16#11#),
      3376 => to_slv(opcode_type, 16#0A#),
      3377 => to_slv(opcode_type, 16#07#),
      3378 => to_slv(opcode_type, 16#0B#),
      3379 => to_slv(opcode_type, 16#0E#),
      3380 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#09#),
      3393 => to_slv(opcode_type, 16#01#),
      3394 => to_slv(opcode_type, 16#04#),
      3395 => to_slv(opcode_type, 16#05#),
      3396 => to_slv(opcode_type, 16#0F#),
      3397 => to_slv(opcode_type, 16#09#),
      3398 => to_slv(opcode_type, 16#06#),
      3399 => to_slv(opcode_type, 16#06#),
      3400 => to_slv(opcode_type, 16#0C#),
      3401 => to_slv(opcode_type, 16#0D#),
      3402 => to_slv(opcode_type, 16#06#),
      3403 => to_slv(opcode_type, 16#0E#),
      3404 => to_slv(opcode_type, 16#DE#),
      3405 => to_slv(opcode_type, 16#06#),
      3406 => to_slv(opcode_type, 16#09#),
      3407 => to_slv(opcode_type, 16#0A#),
      3408 => to_slv(opcode_type, 16#10#),
      3409 => to_slv(opcode_type, 16#06#),
      3410 => to_slv(opcode_type, 16#0F#),
      3411 => to_slv(opcode_type, 16#0D#),
      3412 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#06#),
      3425 => to_slv(opcode_type, 16#07#),
      3426 => to_slv(opcode_type, 16#07#),
      3427 => to_slv(opcode_type, 16#09#),
      3428 => to_slv(opcode_type, 16#0E#),
      3429 => to_slv(opcode_type, 16#10#),
      3430 => to_slv(opcode_type, 16#04#),
      3431 => to_slv(opcode_type, 16#0C#),
      3432 => to_slv(opcode_type, 16#05#),
      3433 => to_slv(opcode_type, 16#06#),
      3434 => to_slv(opcode_type, 16#0D#),
      3435 => to_slv(opcode_type, 16#11#),
      3436 => to_slv(opcode_type, 16#04#),
      3437 => to_slv(opcode_type, 16#09#),
      3438 => to_slv(opcode_type, 16#08#),
      3439 => to_slv(opcode_type, 16#0D#),
      3440 => to_slv(opcode_type, 16#11#),
      3441 => to_slv(opcode_type, 16#08#),
      3442 => to_slv(opcode_type, 16#0B#),
      3443 => to_slv(opcode_type, 16#0B#),
      3444 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#07#),
      3457 => to_slv(opcode_type, 16#05#),
      3458 => to_slv(opcode_type, 16#07#),
      3459 => to_slv(opcode_type, 16#05#),
      3460 => to_slv(opcode_type, 16#0A#),
      3461 => to_slv(opcode_type, 16#05#),
      3462 => to_slv(opcode_type, 16#10#),
      3463 => to_slv(opcode_type, 16#09#),
      3464 => to_slv(opcode_type, 16#09#),
      3465 => to_slv(opcode_type, 16#07#),
      3466 => to_slv(opcode_type, 16#0B#),
      3467 => to_slv(opcode_type, 16#0C#),
      3468 => to_slv(opcode_type, 16#01#),
      3469 => to_slv(opcode_type, 16#10#),
      3470 => to_slv(opcode_type, 16#07#),
      3471 => to_slv(opcode_type, 16#02#),
      3472 => to_slv(opcode_type, 16#29#),
      3473 => to_slv(opcode_type, 16#07#),
      3474 => to_slv(opcode_type, 16#0B#),
      3475 => to_slv(opcode_type, 16#10#),
      3476 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#07#),
      3489 => to_slv(opcode_type, 16#04#),
      3490 => to_slv(opcode_type, 16#03#),
      3491 => to_slv(opcode_type, 16#08#),
      3492 => to_slv(opcode_type, 16#11#),
      3493 => to_slv(opcode_type, 16#0C#),
      3494 => to_slv(opcode_type, 16#07#),
      3495 => to_slv(opcode_type, 16#06#),
      3496 => to_slv(opcode_type, 16#08#),
      3497 => to_slv(opcode_type, 16#0B#),
      3498 => to_slv(opcode_type, 16#0D#),
      3499 => to_slv(opcode_type, 16#04#),
      3500 => to_slv(opcode_type, 16#0A#),
      3501 => to_slv(opcode_type, 16#09#),
      3502 => to_slv(opcode_type, 16#07#),
      3503 => to_slv(opcode_type, 16#11#),
      3504 => to_slv(opcode_type, 16#11#),
      3505 => to_slv(opcode_type, 16#06#),
      3506 => to_slv(opcode_type, 16#0D#),
      3507 => to_slv(opcode_type, 16#10#),
      3508 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#07#),
      3521 => to_slv(opcode_type, 16#06#),
      3522 => to_slv(opcode_type, 16#07#),
      3523 => to_slv(opcode_type, 16#08#),
      3524 => to_slv(opcode_type, 16#0E#),
      3525 => to_slv(opcode_type, 16#0F#),
      3526 => to_slv(opcode_type, 16#02#),
      3527 => to_slv(opcode_type, 16#0F#),
      3528 => to_slv(opcode_type, 16#09#),
      3529 => to_slv(opcode_type, 16#02#),
      3530 => to_slv(opcode_type, 16#0C#),
      3531 => to_slv(opcode_type, 16#03#),
      3532 => to_slv(opcode_type, 16#0D#),
      3533 => to_slv(opcode_type, 16#07#),
      3534 => to_slv(opcode_type, 16#04#),
      3535 => to_slv(opcode_type, 16#08#),
      3536 => to_slv(opcode_type, 16#0D#),
      3537 => to_slv(opcode_type, 16#0B#),
      3538 => to_slv(opcode_type, 16#02#),
      3539 => to_slv(opcode_type, 16#0F#),
      3540 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#06#),
      3553 => to_slv(opcode_type, 16#03#),
      3554 => to_slv(opcode_type, 16#07#),
      3555 => to_slv(opcode_type, 16#04#),
      3556 => to_slv(opcode_type, 16#88#),
      3557 => to_slv(opcode_type, 16#01#),
      3558 => to_slv(opcode_type, 16#0F#),
      3559 => to_slv(opcode_type, 16#09#),
      3560 => to_slv(opcode_type, 16#07#),
      3561 => to_slv(opcode_type, 16#04#),
      3562 => to_slv(opcode_type, 16#10#),
      3563 => to_slv(opcode_type, 16#05#),
      3564 => to_slv(opcode_type, 16#11#),
      3565 => to_slv(opcode_type, 16#06#),
      3566 => to_slv(opcode_type, 16#06#),
      3567 => to_slv(opcode_type, 16#CD#),
      3568 => to_slv(opcode_type, 16#10#),
      3569 => to_slv(opcode_type, 16#09#),
      3570 => to_slv(opcode_type, 16#0E#),
      3571 => to_slv(opcode_type, 16#0B#),
      3572 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#08#),
      3585 => to_slv(opcode_type, 16#01#),
      3586 => to_slv(opcode_type, 16#08#),
      3587 => to_slv(opcode_type, 16#06#),
      3588 => to_slv(opcode_type, 16#0A#),
      3589 => to_slv(opcode_type, 16#10#),
      3590 => to_slv(opcode_type, 16#01#),
      3591 => to_slv(opcode_type, 16#11#),
      3592 => to_slv(opcode_type, 16#09#),
      3593 => to_slv(opcode_type, 16#04#),
      3594 => to_slv(opcode_type, 16#09#),
      3595 => to_slv(opcode_type, 16#11#),
      3596 => to_slv(opcode_type, 16#0E#),
      3597 => to_slv(opcode_type, 16#07#),
      3598 => to_slv(opcode_type, 16#09#),
      3599 => to_slv(opcode_type, 16#0C#),
      3600 => to_slv(opcode_type, 16#97#),
      3601 => to_slv(opcode_type, 16#09#),
      3602 => to_slv(opcode_type, 16#0B#),
      3603 => to_slv(opcode_type, 16#F8#),
      3604 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#09#),
      3617 => to_slv(opcode_type, 16#03#),
      3618 => to_slv(opcode_type, 16#08#),
      3619 => to_slv(opcode_type, 16#04#),
      3620 => to_slv(opcode_type, 16#C5#),
      3621 => to_slv(opcode_type, 16#07#),
      3622 => to_slv(opcode_type, 16#A4#),
      3623 => to_slv(opcode_type, 16#0D#),
      3624 => to_slv(opcode_type, 16#06#),
      3625 => to_slv(opcode_type, 16#04#),
      3626 => to_slv(opcode_type, 16#06#),
      3627 => to_slv(opcode_type, 16#0B#),
      3628 => to_slv(opcode_type, 16#11#),
      3629 => to_slv(opcode_type, 16#08#),
      3630 => to_slv(opcode_type, 16#06#),
      3631 => to_slv(opcode_type, 16#AB#),
      3632 => to_slv(opcode_type, 16#0F#),
      3633 => to_slv(opcode_type, 16#09#),
      3634 => to_slv(opcode_type, 16#0A#),
      3635 => to_slv(opcode_type, 16#0D#),
      3636 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#06#),
      3649 => to_slv(opcode_type, 16#03#),
      3650 => to_slv(opcode_type, 16#06#),
      3651 => to_slv(opcode_type, 16#01#),
      3652 => to_slv(opcode_type, 16#0B#),
      3653 => to_slv(opcode_type, 16#04#),
      3654 => to_slv(opcode_type, 16#0D#),
      3655 => to_slv(opcode_type, 16#08#),
      3656 => to_slv(opcode_type, 16#07#),
      3657 => to_slv(opcode_type, 16#06#),
      3658 => to_slv(opcode_type, 16#0C#),
      3659 => to_slv(opcode_type, 16#0B#),
      3660 => to_slv(opcode_type, 16#04#),
      3661 => to_slv(opcode_type, 16#11#),
      3662 => to_slv(opcode_type, 16#07#),
      3663 => to_slv(opcode_type, 16#07#),
      3664 => to_slv(opcode_type, 16#0E#),
      3665 => to_slv(opcode_type, 16#0B#),
      3666 => to_slv(opcode_type, 16#01#),
      3667 => to_slv(opcode_type, 16#0B#),
      3668 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#08#),
      3681 => to_slv(opcode_type, 16#06#),
      3682 => to_slv(opcode_type, 16#02#),
      3683 => to_slv(opcode_type, 16#05#),
      3684 => to_slv(opcode_type, 16#64#),
      3685 => to_slv(opcode_type, 16#09#),
      3686 => to_slv(opcode_type, 16#07#),
      3687 => to_slv(opcode_type, 16#0D#),
      3688 => to_slv(opcode_type, 16#0E#),
      3689 => to_slv(opcode_type, 16#09#),
      3690 => to_slv(opcode_type, 16#0F#),
      3691 => to_slv(opcode_type, 16#26#),
      3692 => to_slv(opcode_type, 16#09#),
      3693 => to_slv(opcode_type, 16#01#),
      3694 => to_slv(opcode_type, 16#02#),
      3695 => to_slv(opcode_type, 16#10#),
      3696 => to_slv(opcode_type, 16#03#),
      3697 => to_slv(opcode_type, 16#07#),
      3698 => to_slv(opcode_type, 16#96#),
      3699 => to_slv(opcode_type, 16#11#),
      3700 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#08#),
      3713 => to_slv(opcode_type, 16#05#),
      3714 => to_slv(opcode_type, 16#01#),
      3715 => to_slv(opcode_type, 16#08#),
      3716 => to_slv(opcode_type, 16#0F#),
      3717 => to_slv(opcode_type, 16#0D#),
      3718 => to_slv(opcode_type, 16#09#),
      3719 => to_slv(opcode_type, 16#06#),
      3720 => to_slv(opcode_type, 16#01#),
      3721 => to_slv(opcode_type, 16#0F#),
      3722 => to_slv(opcode_type, 16#06#),
      3723 => to_slv(opcode_type, 16#11#),
      3724 => to_slv(opcode_type, 16#0B#),
      3725 => to_slv(opcode_type, 16#09#),
      3726 => to_slv(opcode_type, 16#07#),
      3727 => to_slv(opcode_type, 16#0A#),
      3728 => to_slv(opcode_type, 16#0C#),
      3729 => to_slv(opcode_type, 16#07#),
      3730 => to_slv(opcode_type, 16#0D#),
      3731 => to_slv(opcode_type, 16#0D#),
      3732 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#08#),
      3745 => to_slv(opcode_type, 16#08#),
      3746 => to_slv(opcode_type, 16#05#),
      3747 => to_slv(opcode_type, 16#09#),
      3748 => to_slv(opcode_type, 16#E4#),
      3749 => to_slv(opcode_type, 16#0B#),
      3750 => to_slv(opcode_type, 16#02#),
      3751 => to_slv(opcode_type, 16#03#),
      3752 => to_slv(opcode_type, 16#0F#),
      3753 => to_slv(opcode_type, 16#06#),
      3754 => to_slv(opcode_type, 16#01#),
      3755 => to_slv(opcode_type, 16#05#),
      3756 => to_slv(opcode_type, 16#0C#),
      3757 => to_slv(opcode_type, 16#08#),
      3758 => to_slv(opcode_type, 16#07#),
      3759 => to_slv(opcode_type, 16#A3#),
      3760 => to_slv(opcode_type, 16#0F#),
      3761 => to_slv(opcode_type, 16#09#),
      3762 => to_slv(opcode_type, 16#0A#),
      3763 => to_slv(opcode_type, 16#99#),
      3764 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#08#),
      3777 => to_slv(opcode_type, 16#06#),
      3778 => to_slv(opcode_type, 16#08#),
      3779 => to_slv(opcode_type, 16#03#),
      3780 => to_slv(opcode_type, 16#0B#),
      3781 => to_slv(opcode_type, 16#05#),
      3782 => to_slv(opcode_type, 16#0B#),
      3783 => to_slv(opcode_type, 16#08#),
      3784 => to_slv(opcode_type, 16#07#),
      3785 => to_slv(opcode_type, 16#0A#),
      3786 => to_slv(opcode_type, 16#0E#),
      3787 => to_slv(opcode_type, 16#01#),
      3788 => to_slv(opcode_type, 16#11#),
      3789 => to_slv(opcode_type, 16#08#),
      3790 => to_slv(opcode_type, 16#08#),
      3791 => to_slv(opcode_type, 16#03#),
      3792 => to_slv(opcode_type, 16#11#),
      3793 => to_slv(opcode_type, 16#02#),
      3794 => to_slv(opcode_type, 16#0A#),
      3795 => to_slv(opcode_type, 16#0B#),
      3796 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#09#),
      3809 => to_slv(opcode_type, 16#05#),
      3810 => to_slv(opcode_type, 16#07#),
      3811 => to_slv(opcode_type, 16#03#),
      3812 => to_slv(opcode_type, 16#0B#),
      3813 => to_slv(opcode_type, 16#08#),
      3814 => to_slv(opcode_type, 16#0C#),
      3815 => to_slv(opcode_type, 16#11#),
      3816 => to_slv(opcode_type, 16#06#),
      3817 => to_slv(opcode_type, 16#08#),
      3818 => to_slv(opcode_type, 16#02#),
      3819 => to_slv(opcode_type, 16#0A#),
      3820 => to_slv(opcode_type, 16#06#),
      3821 => to_slv(opcode_type, 16#0F#),
      3822 => to_slv(opcode_type, 16#0E#),
      3823 => to_slv(opcode_type, 16#08#),
      3824 => to_slv(opcode_type, 16#07#),
      3825 => to_slv(opcode_type, 16#0C#),
      3826 => to_slv(opcode_type, 16#0A#),
      3827 => to_slv(opcode_type, 16#0E#),
      3828 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#07#),
      3841 => to_slv(opcode_type, 16#06#),
      3842 => to_slv(opcode_type, 16#04#),
      3843 => to_slv(opcode_type, 16#09#),
      3844 => to_slv(opcode_type, 16#0B#),
      3845 => to_slv(opcode_type, 16#0B#),
      3846 => to_slv(opcode_type, 16#04#),
      3847 => to_slv(opcode_type, 16#07#),
      3848 => to_slv(opcode_type, 16#0E#),
      3849 => to_slv(opcode_type, 16#0C#),
      3850 => to_slv(opcode_type, 16#08#),
      3851 => to_slv(opcode_type, 16#06#),
      3852 => to_slv(opcode_type, 16#07#),
      3853 => to_slv(opcode_type, 16#0A#),
      3854 => to_slv(opcode_type, 16#0B#),
      3855 => to_slv(opcode_type, 16#09#),
      3856 => to_slv(opcode_type, 16#0F#),
      3857 => to_slv(opcode_type, 16#E6#),
      3858 => to_slv(opcode_type, 16#01#),
      3859 => to_slv(opcode_type, 16#0D#),
      3860 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#09#),
      3873 => to_slv(opcode_type, 16#06#),
      3874 => to_slv(opcode_type, 16#05#),
      3875 => to_slv(opcode_type, 16#09#),
      3876 => to_slv(opcode_type, 16#0D#),
      3877 => to_slv(opcode_type, 16#0D#),
      3878 => to_slv(opcode_type, 16#07#),
      3879 => to_slv(opcode_type, 16#07#),
      3880 => to_slv(opcode_type, 16#0D#),
      3881 => to_slv(opcode_type, 16#0D#),
      3882 => to_slv(opcode_type, 16#04#),
      3883 => to_slv(opcode_type, 16#0A#),
      3884 => to_slv(opcode_type, 16#03#),
      3885 => to_slv(opcode_type, 16#09#),
      3886 => to_slv(opcode_type, 16#08#),
      3887 => to_slv(opcode_type, 16#10#),
      3888 => to_slv(opcode_type, 16#0B#),
      3889 => to_slv(opcode_type, 16#08#),
      3890 => to_slv(opcode_type, 16#0F#),
      3891 => to_slv(opcode_type, 16#0F#),
      3892 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#09#),
      3905 => to_slv(opcode_type, 16#09#),
      3906 => to_slv(opcode_type, 16#06#),
      3907 => to_slv(opcode_type, 16#03#),
      3908 => to_slv(opcode_type, 16#11#),
      3909 => to_slv(opcode_type, 16#03#),
      3910 => to_slv(opcode_type, 16#0E#),
      3911 => to_slv(opcode_type, 16#03#),
      3912 => to_slv(opcode_type, 16#03#),
      3913 => to_slv(opcode_type, 16#40#),
      3914 => to_slv(opcode_type, 16#06#),
      3915 => to_slv(opcode_type, 16#04#),
      3916 => to_slv(opcode_type, 16#05#),
      3917 => to_slv(opcode_type, 16#0A#),
      3918 => to_slv(opcode_type, 16#06#),
      3919 => to_slv(opcode_type, 16#02#),
      3920 => to_slv(opcode_type, 16#0A#),
      3921 => to_slv(opcode_type, 16#09#),
      3922 => to_slv(opcode_type, 16#0E#),
      3923 => to_slv(opcode_type, 16#0C#),
      3924 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#06#),
      3937 => to_slv(opcode_type, 16#04#),
      3938 => to_slv(opcode_type, 16#03#),
      3939 => to_slv(opcode_type, 16#09#),
      3940 => to_slv(opcode_type, 16#10#),
      3941 => to_slv(opcode_type, 16#0C#),
      3942 => to_slv(opcode_type, 16#09#),
      3943 => to_slv(opcode_type, 16#06#),
      3944 => to_slv(opcode_type, 16#05#),
      3945 => to_slv(opcode_type, 16#10#),
      3946 => to_slv(opcode_type, 16#09#),
      3947 => to_slv(opcode_type, 16#0D#),
      3948 => to_slv(opcode_type, 16#0E#),
      3949 => to_slv(opcode_type, 16#08#),
      3950 => to_slv(opcode_type, 16#06#),
      3951 => to_slv(opcode_type, 16#0C#),
      3952 => to_slv(opcode_type, 16#0D#),
      3953 => to_slv(opcode_type, 16#09#),
      3954 => to_slv(opcode_type, 16#11#),
      3955 => to_slv(opcode_type, 16#0A#),
      3956 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#06#),
      3969 => to_slv(opcode_type, 16#07#),
      3970 => to_slv(opcode_type, 16#05#),
      3971 => to_slv(opcode_type, 16#09#),
      3972 => to_slv(opcode_type, 16#0F#),
      3973 => to_slv(opcode_type, 16#0B#),
      3974 => to_slv(opcode_type, 16#09#),
      3975 => to_slv(opcode_type, 16#09#),
      3976 => to_slv(opcode_type, 16#0B#),
      3977 => to_slv(opcode_type, 16#11#),
      3978 => to_slv(opcode_type, 16#05#),
      3979 => to_slv(opcode_type, 16#0E#),
      3980 => to_slv(opcode_type, 16#03#),
      3981 => to_slv(opcode_type, 16#08#),
      3982 => to_slv(opcode_type, 16#08#),
      3983 => to_slv(opcode_type, 16#0F#),
      3984 => to_slv(opcode_type, 16#11#),
      3985 => to_slv(opcode_type, 16#09#),
      3986 => to_slv(opcode_type, 16#11#),
      3987 => to_slv(opcode_type, 16#10#),
      3988 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#07#),
      4001 => to_slv(opcode_type, 16#01#),
      4002 => to_slv(opcode_type, 16#07#),
      4003 => to_slv(opcode_type, 16#01#),
      4004 => to_slv(opcode_type, 16#0A#),
      4005 => to_slv(opcode_type, 16#05#),
      4006 => to_slv(opcode_type, 16#10#),
      4007 => to_slv(opcode_type, 16#09#),
      4008 => to_slv(opcode_type, 16#09#),
      4009 => to_slv(opcode_type, 16#03#),
      4010 => to_slv(opcode_type, 16#11#),
      4011 => to_slv(opcode_type, 16#05#),
      4012 => to_slv(opcode_type, 16#0A#),
      4013 => to_slv(opcode_type, 16#09#),
      4014 => to_slv(opcode_type, 16#09#),
      4015 => to_slv(opcode_type, 16#0B#),
      4016 => to_slv(opcode_type, 16#0D#),
      4017 => to_slv(opcode_type, 16#08#),
      4018 => to_slv(opcode_type, 16#0F#),
      4019 => to_slv(opcode_type, 16#10#),
      4020 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#09#),
      4033 => to_slv(opcode_type, 16#01#),
      4034 => to_slv(opcode_type, 16#06#),
      4035 => to_slv(opcode_type, 16#04#),
      4036 => to_slv(opcode_type, 16#BF#),
      4037 => to_slv(opcode_type, 16#01#),
      4038 => to_slv(opcode_type, 16#0A#),
      4039 => to_slv(opcode_type, 16#06#),
      4040 => to_slv(opcode_type, 16#09#),
      4041 => to_slv(opcode_type, 16#09#),
      4042 => to_slv(opcode_type, 16#0B#),
      4043 => to_slv(opcode_type, 16#0B#),
      4044 => to_slv(opcode_type, 16#01#),
      4045 => to_slv(opcode_type, 16#0B#),
      4046 => to_slv(opcode_type, 16#08#),
      4047 => to_slv(opcode_type, 16#09#),
      4048 => to_slv(opcode_type, 16#0A#),
      4049 => to_slv(opcode_type, 16#11#),
      4050 => to_slv(opcode_type, 16#04#),
      4051 => to_slv(opcode_type, 16#10#),
      4052 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#04#),
      4066 => to_slv(opcode_type, 16#01#),
      4067 => to_slv(opcode_type, 16#04#),
      4068 => to_slv(opcode_type, 16#0D#),
      4069 => to_slv(opcode_type, 16#06#),
      4070 => to_slv(opcode_type, 16#09#),
      4071 => to_slv(opcode_type, 16#09#),
      4072 => to_slv(opcode_type, 16#0E#),
      4073 => to_slv(opcode_type, 16#0C#),
      4074 => to_slv(opcode_type, 16#09#),
      4075 => to_slv(opcode_type, 16#0C#),
      4076 => to_slv(opcode_type, 16#11#),
      4077 => to_slv(opcode_type, 16#07#),
      4078 => to_slv(opcode_type, 16#09#),
      4079 => to_slv(opcode_type, 16#FC#),
      4080 => to_slv(opcode_type, 16#0C#),
      4081 => to_slv(opcode_type, 16#06#),
      4082 => to_slv(opcode_type, 16#0F#),
      4083 => to_slv(opcode_type, 16#0C#),
      4084 to 4095 => (others => '0')
  ),

    -- Bin `21`...
    20 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#09#),
      1 => to_slv(opcode_type, 16#05#),
      2 => to_slv(opcode_type, 16#08#),
      3 => to_slv(opcode_type, 16#08#),
      4 => to_slv(opcode_type, 16#0F#),
      5 => to_slv(opcode_type, 16#0F#),
      6 => to_slv(opcode_type, 16#05#),
      7 => to_slv(opcode_type, 16#0F#),
      8 => to_slv(opcode_type, 16#09#),
      9 => to_slv(opcode_type, 16#06#),
      10 => to_slv(opcode_type, 16#05#),
      11 => to_slv(opcode_type, 16#10#),
      12 => to_slv(opcode_type, 16#08#),
      13 => to_slv(opcode_type, 16#0A#),
      14 => to_slv(opcode_type, 16#0C#),
      15 => to_slv(opcode_type, 16#06#),
      16 => to_slv(opcode_type, 16#06#),
      17 => to_slv(opcode_type, 16#0F#),
      18 => to_slv(opcode_type, 16#0E#),
      19 => to_slv(opcode_type, 16#02#),
      20 => to_slv(opcode_type, 16#0C#),
      21 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#09#),
      33 => to_slv(opcode_type, 16#01#),
      34 => to_slv(opcode_type, 16#09#),
      35 => to_slv(opcode_type, 16#04#),
      36 => to_slv(opcode_type, 16#0B#),
      37 => to_slv(opcode_type, 16#02#),
      38 => to_slv(opcode_type, 16#10#),
      39 => to_slv(opcode_type, 16#06#),
      40 => to_slv(opcode_type, 16#08#),
      41 => to_slv(opcode_type, 16#02#),
      42 => to_slv(opcode_type, 16#0F#),
      43 => to_slv(opcode_type, 16#07#),
      44 => to_slv(opcode_type, 16#11#),
      45 => to_slv(opcode_type, 16#1F#),
      46 => to_slv(opcode_type, 16#06#),
      47 => to_slv(opcode_type, 16#06#),
      48 => to_slv(opcode_type, 16#0C#),
      49 => to_slv(opcode_type, 16#0C#),
      50 => to_slv(opcode_type, 16#06#),
      51 => to_slv(opcode_type, 16#0F#),
      52 => to_slv(opcode_type, 16#0F#),
      53 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#08#),
      65 => to_slv(opcode_type, 16#06#),
      66 => to_slv(opcode_type, 16#01#),
      67 => to_slv(opcode_type, 16#02#),
      68 => to_slv(opcode_type, 16#0C#),
      69 => to_slv(opcode_type, 16#04#),
      70 => to_slv(opcode_type, 16#07#),
      71 => to_slv(opcode_type, 16#0F#),
      72 => to_slv(opcode_type, 16#0C#),
      73 => to_slv(opcode_type, 16#07#),
      74 => to_slv(opcode_type, 16#07#),
      75 => to_slv(opcode_type, 16#06#),
      76 => to_slv(opcode_type, 16#10#),
      77 => to_slv(opcode_type, 16#0F#),
      78 => to_slv(opcode_type, 16#05#),
      79 => to_slv(opcode_type, 16#10#),
      80 => to_slv(opcode_type, 16#07#),
      81 => to_slv(opcode_type, 16#07#),
      82 => to_slv(opcode_type, 16#0D#),
      83 => to_slv(opcode_type, 16#11#),
      84 => to_slv(opcode_type, 16#0E#),
      85 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#09#),
      97 => to_slv(opcode_type, 16#09#),
      98 => to_slv(opcode_type, 16#02#),
      99 => to_slv(opcode_type, 16#08#),
      100 => to_slv(opcode_type, 16#0A#),
      101 => to_slv(opcode_type, 16#0F#),
      102 => to_slv(opcode_type, 16#06#),
      103 => to_slv(opcode_type, 16#08#),
      104 => to_slv(opcode_type, 16#11#),
      105 => to_slv(opcode_type, 16#0C#),
      106 => to_slv(opcode_type, 16#03#),
      107 => to_slv(opcode_type, 16#0F#),
      108 => to_slv(opcode_type, 16#07#),
      109 => to_slv(opcode_type, 16#07#),
      110 => to_slv(opcode_type, 16#02#),
      111 => to_slv(opcode_type, 16#0C#),
      112 => to_slv(opcode_type, 16#03#),
      113 => to_slv(opcode_type, 16#11#),
      114 => to_slv(opcode_type, 16#05#),
      115 => to_slv(opcode_type, 16#05#),
      116 => to_slv(opcode_type, 16#E4#),
      117 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#06#),
      129 => to_slv(opcode_type, 16#02#),
      130 => to_slv(opcode_type, 16#03#),
      131 => to_slv(opcode_type, 16#06#),
      132 => to_slv(opcode_type, 16#0C#),
      133 => to_slv(opcode_type, 16#10#),
      134 => to_slv(opcode_type, 16#06#),
      135 => to_slv(opcode_type, 16#08#),
      136 => to_slv(opcode_type, 16#08#),
      137 => to_slv(opcode_type, 16#0E#),
      138 => to_slv(opcode_type, 16#11#),
      139 => to_slv(opcode_type, 16#06#),
      140 => to_slv(opcode_type, 16#0F#),
      141 => to_slv(opcode_type, 16#11#),
      142 => to_slv(opcode_type, 16#08#),
      143 => to_slv(opcode_type, 16#06#),
      144 => to_slv(opcode_type, 16#10#),
      145 => to_slv(opcode_type, 16#0F#),
      146 => to_slv(opcode_type, 16#07#),
      147 => to_slv(opcode_type, 16#0C#),
      148 => to_slv(opcode_type, 16#5B#),
      149 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#09#),
      161 => to_slv(opcode_type, 16#08#),
      162 => to_slv(opcode_type, 16#08#),
      163 => to_slv(opcode_type, 16#09#),
      164 => to_slv(opcode_type, 16#0C#),
      165 => to_slv(opcode_type, 16#AF#),
      166 => to_slv(opcode_type, 16#05#),
      167 => to_slv(opcode_type, 16#11#),
      168 => to_slv(opcode_type, 16#09#),
      169 => to_slv(opcode_type, 16#05#),
      170 => to_slv(opcode_type, 16#0E#),
      171 => to_slv(opcode_type, 16#06#),
      172 => to_slv(opcode_type, 16#D6#),
      173 => to_slv(opcode_type, 16#0D#),
      174 => to_slv(opcode_type, 16#06#),
      175 => to_slv(opcode_type, 16#09#),
      176 => to_slv(opcode_type, 16#06#),
      177 => to_slv(opcode_type, 16#84#),
      178 => to_slv(opcode_type, 16#0D#),
      179 => to_slv(opcode_type, 16#0D#),
      180 => to_slv(opcode_type, 16#10#),
      181 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#07#),
      193 => to_slv(opcode_type, 16#08#),
      194 => to_slv(opcode_type, 16#07#),
      195 => to_slv(opcode_type, 16#04#),
      196 => to_slv(opcode_type, 16#0C#),
      197 => to_slv(opcode_type, 16#07#),
      198 => to_slv(opcode_type, 16#0D#),
      199 => to_slv(opcode_type, 16#10#),
      200 => to_slv(opcode_type, 16#08#),
      201 => to_slv(opcode_type, 16#02#),
      202 => to_slv(opcode_type, 16#11#),
      203 => to_slv(opcode_type, 16#05#),
      204 => to_slv(opcode_type, 16#10#),
      205 => to_slv(opcode_type, 16#03#),
      206 => to_slv(opcode_type, 16#06#),
      207 => to_slv(opcode_type, 16#07#),
      208 => to_slv(opcode_type, 16#0F#),
      209 => to_slv(opcode_type, 16#0B#),
      210 => to_slv(opcode_type, 16#06#),
      211 => to_slv(opcode_type, 16#0B#),
      212 => to_slv(opcode_type, 16#1D#),
      213 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#09#),
      225 => to_slv(opcode_type, 16#05#),
      226 => to_slv(opcode_type, 16#03#),
      227 => to_slv(opcode_type, 16#08#),
      228 => to_slv(opcode_type, 16#11#),
      229 => to_slv(opcode_type, 16#0B#),
      230 => to_slv(opcode_type, 16#08#),
      231 => to_slv(opcode_type, 16#09#),
      232 => to_slv(opcode_type, 16#07#),
      233 => to_slv(opcode_type, 16#B5#),
      234 => to_slv(opcode_type, 16#10#),
      235 => to_slv(opcode_type, 16#06#),
      236 => to_slv(opcode_type, 16#0A#),
      237 => to_slv(opcode_type, 16#0C#),
      238 => to_slv(opcode_type, 16#09#),
      239 => to_slv(opcode_type, 16#06#),
      240 => to_slv(opcode_type, 16#11#),
      241 => to_slv(opcode_type, 16#0F#),
      242 => to_slv(opcode_type, 16#07#),
      243 => to_slv(opcode_type, 16#0C#),
      244 => to_slv(opcode_type, 16#0C#),
      245 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#08#),
      257 => to_slv(opcode_type, 16#09#),
      258 => to_slv(opcode_type, 16#08#),
      259 => to_slv(opcode_type, 16#06#),
      260 => to_slv(opcode_type, 16#0C#),
      261 => to_slv(opcode_type, 16#0B#),
      262 => to_slv(opcode_type, 16#04#),
      263 => to_slv(opcode_type, 16#0F#),
      264 => to_slv(opcode_type, 16#03#),
      265 => to_slv(opcode_type, 16#09#),
      266 => to_slv(opcode_type, 16#0B#),
      267 => to_slv(opcode_type, 16#0B#),
      268 => to_slv(opcode_type, 16#07#),
      269 => to_slv(opcode_type, 16#06#),
      270 => to_slv(opcode_type, 16#09#),
      271 => to_slv(opcode_type, 16#31#),
      272 => to_slv(opcode_type, 16#0B#),
      273 => to_slv(opcode_type, 16#08#),
      274 => to_slv(opcode_type, 16#0F#),
      275 => to_slv(opcode_type, 16#0C#),
      276 => to_slv(opcode_type, 16#0D#),
      277 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#09#),
      290 => to_slv(opcode_type, 16#01#),
      291 => to_slv(opcode_type, 16#02#),
      292 => to_slv(opcode_type, 16#0C#),
      293 => to_slv(opcode_type, 16#01#),
      294 => to_slv(opcode_type, 16#02#),
      295 => to_slv(opcode_type, 16#0F#),
      296 => to_slv(opcode_type, 16#07#),
      297 => to_slv(opcode_type, 16#09#),
      298 => to_slv(opcode_type, 16#07#),
      299 => to_slv(opcode_type, 16#0E#),
      300 => to_slv(opcode_type, 16#0C#),
      301 => to_slv(opcode_type, 16#02#),
      302 => to_slv(opcode_type, 16#11#),
      303 => to_slv(opcode_type, 16#08#),
      304 => to_slv(opcode_type, 16#01#),
      305 => to_slv(opcode_type, 16#D4#),
      306 => to_slv(opcode_type, 16#08#),
      307 => to_slv(opcode_type, 16#0E#),
      308 => to_slv(opcode_type, 16#11#),
      309 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#06#),
      321 => to_slv(opcode_type, 16#08#),
      322 => to_slv(opcode_type, 16#09#),
      323 => to_slv(opcode_type, 16#07#),
      324 => to_slv(opcode_type, 16#0F#),
      325 => to_slv(opcode_type, 16#10#),
      326 => to_slv(opcode_type, 16#06#),
      327 => to_slv(opcode_type, 16#0D#),
      328 => to_slv(opcode_type, 16#10#),
      329 => to_slv(opcode_type, 16#02#),
      330 => to_slv(opcode_type, 16#04#),
      331 => to_slv(opcode_type, 16#0D#),
      332 => to_slv(opcode_type, 16#07#),
      333 => to_slv(opcode_type, 16#05#),
      334 => to_slv(opcode_type, 16#03#),
      335 => to_slv(opcode_type, 16#0C#),
      336 => to_slv(opcode_type, 16#07#),
      337 => to_slv(opcode_type, 16#05#),
      338 => to_slv(opcode_type, 16#0A#),
      339 => to_slv(opcode_type, 16#03#),
      340 => to_slv(opcode_type, 16#11#),
      341 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#06#),
      353 => to_slv(opcode_type, 16#05#),
      354 => to_slv(opcode_type, 16#05#),
      355 => to_slv(opcode_type, 16#08#),
      356 => to_slv(opcode_type, 16#10#),
      357 => to_slv(opcode_type, 16#0B#),
      358 => to_slv(opcode_type, 16#08#),
      359 => to_slv(opcode_type, 16#07#),
      360 => to_slv(opcode_type, 16#08#),
      361 => to_slv(opcode_type, 16#0A#),
      362 => to_slv(opcode_type, 16#0C#),
      363 => to_slv(opcode_type, 16#07#),
      364 => to_slv(opcode_type, 16#0E#),
      365 => to_slv(opcode_type, 16#65#),
      366 => to_slv(opcode_type, 16#06#),
      367 => to_slv(opcode_type, 16#06#),
      368 => to_slv(opcode_type, 16#0E#),
      369 => to_slv(opcode_type, 16#0E#),
      370 => to_slv(opcode_type, 16#08#),
      371 => to_slv(opcode_type, 16#0E#),
      372 => to_slv(opcode_type, 16#0F#),
      373 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#06#),
      385 => to_slv(opcode_type, 16#04#),
      386 => to_slv(opcode_type, 16#04#),
      387 => to_slv(opcode_type, 16#06#),
      388 => to_slv(opcode_type, 16#0B#),
      389 => to_slv(opcode_type, 16#11#),
      390 => to_slv(opcode_type, 16#06#),
      391 => to_slv(opcode_type, 16#08#),
      392 => to_slv(opcode_type, 16#09#),
      393 => to_slv(opcode_type, 16#0E#),
      394 => to_slv(opcode_type, 16#0E#),
      395 => to_slv(opcode_type, 16#07#),
      396 => to_slv(opcode_type, 16#10#),
      397 => to_slv(opcode_type, 16#11#),
      398 => to_slv(opcode_type, 16#08#),
      399 => to_slv(opcode_type, 16#08#),
      400 => to_slv(opcode_type, 16#10#),
      401 => to_slv(opcode_type, 16#0A#),
      402 => to_slv(opcode_type, 16#07#),
      403 => to_slv(opcode_type, 16#0E#),
      404 => to_slv(opcode_type, 16#10#),
      405 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#07#),
      417 => to_slv(opcode_type, 16#07#),
      418 => to_slv(opcode_type, 16#03#),
      419 => to_slv(opcode_type, 16#07#),
      420 => to_slv(opcode_type, 16#11#),
      421 => to_slv(opcode_type, 16#11#),
      422 => to_slv(opcode_type, 16#09#),
      423 => to_slv(opcode_type, 16#06#),
      424 => to_slv(opcode_type, 16#11#),
      425 => to_slv(opcode_type, 16#0F#),
      426 => to_slv(opcode_type, 16#03#),
      427 => to_slv(opcode_type, 16#0B#),
      428 => to_slv(opcode_type, 16#08#),
      429 => to_slv(opcode_type, 16#06#),
      430 => to_slv(opcode_type, 16#02#),
      431 => to_slv(opcode_type, 16#11#),
      432 => to_slv(opcode_type, 16#05#),
      433 => to_slv(opcode_type, 16#0B#),
      434 => to_slv(opcode_type, 16#07#),
      435 => to_slv(opcode_type, 16#10#),
      436 => to_slv(opcode_type, 16#0D#),
      437 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#06#),
      449 => to_slv(opcode_type, 16#03#),
      450 => to_slv(opcode_type, 16#05#),
      451 => to_slv(opcode_type, 16#06#),
      452 => to_slv(opcode_type, 16#0A#),
      453 => to_slv(opcode_type, 16#0B#),
      454 => to_slv(opcode_type, 16#08#),
      455 => to_slv(opcode_type, 16#09#),
      456 => to_slv(opcode_type, 16#06#),
      457 => to_slv(opcode_type, 16#0B#),
      458 => to_slv(opcode_type, 16#10#),
      459 => to_slv(opcode_type, 16#09#),
      460 => to_slv(opcode_type, 16#11#),
      461 => to_slv(opcode_type, 16#0E#),
      462 => to_slv(opcode_type, 16#06#),
      463 => to_slv(opcode_type, 16#07#),
      464 => to_slv(opcode_type, 16#11#),
      465 => to_slv(opcode_type, 16#10#),
      466 => to_slv(opcode_type, 16#06#),
      467 => to_slv(opcode_type, 16#11#),
      468 => to_slv(opcode_type, 16#0C#),
      469 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#08#),
      481 => to_slv(opcode_type, 16#03#),
      482 => to_slv(opcode_type, 16#09#),
      483 => to_slv(opcode_type, 16#02#),
      484 => to_slv(opcode_type, 16#12#),
      485 => to_slv(opcode_type, 16#08#),
      486 => to_slv(opcode_type, 16#B2#),
      487 => to_slv(opcode_type, 16#44#),
      488 => to_slv(opcode_type, 16#09#),
      489 => to_slv(opcode_type, 16#07#),
      490 => to_slv(opcode_type, 16#06#),
      491 => to_slv(opcode_type, 16#0D#),
      492 => to_slv(opcode_type, 16#0E#),
      493 => to_slv(opcode_type, 16#01#),
      494 => to_slv(opcode_type, 16#0B#),
      495 => to_slv(opcode_type, 16#06#),
      496 => to_slv(opcode_type, 16#07#),
      497 => to_slv(opcode_type, 16#0C#),
      498 => to_slv(opcode_type, 16#0D#),
      499 => to_slv(opcode_type, 16#01#),
      500 => to_slv(opcode_type, 16#0A#),
      501 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#07#),
      513 => to_slv(opcode_type, 16#03#),
      514 => to_slv(opcode_type, 16#03#),
      515 => to_slv(opcode_type, 16#06#),
      516 => to_slv(opcode_type, 16#E6#),
      517 => to_slv(opcode_type, 16#DE#),
      518 => to_slv(opcode_type, 16#08#),
      519 => to_slv(opcode_type, 16#06#),
      520 => to_slv(opcode_type, 16#08#),
      521 => to_slv(opcode_type, 16#0E#),
      522 => to_slv(opcode_type, 16#11#),
      523 => to_slv(opcode_type, 16#09#),
      524 => to_slv(opcode_type, 16#B4#),
      525 => to_slv(opcode_type, 16#7D#),
      526 => to_slv(opcode_type, 16#06#),
      527 => to_slv(opcode_type, 16#09#),
      528 => to_slv(opcode_type, 16#0F#),
      529 => to_slv(opcode_type, 16#0E#),
      530 => to_slv(opcode_type, 16#09#),
      531 => to_slv(opcode_type, 16#0C#),
      532 => to_slv(opcode_type, 16#0F#),
      533 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#07#),
      545 => to_slv(opcode_type, 16#04#),
      546 => to_slv(opcode_type, 16#03#),
      547 => to_slv(opcode_type, 16#06#),
      548 => to_slv(opcode_type, 16#0B#),
      549 => to_slv(opcode_type, 16#0C#),
      550 => to_slv(opcode_type, 16#08#),
      551 => to_slv(opcode_type, 16#07#),
      552 => to_slv(opcode_type, 16#06#),
      553 => to_slv(opcode_type, 16#0C#),
      554 => to_slv(opcode_type, 16#0C#),
      555 => to_slv(opcode_type, 16#09#),
      556 => to_slv(opcode_type, 16#0C#),
      557 => to_slv(opcode_type, 16#0D#),
      558 => to_slv(opcode_type, 16#07#),
      559 => to_slv(opcode_type, 16#07#),
      560 => to_slv(opcode_type, 16#0B#),
      561 => to_slv(opcode_type, 16#0B#),
      562 => to_slv(opcode_type, 16#09#),
      563 => to_slv(opcode_type, 16#0D#),
      564 => to_slv(opcode_type, 16#0E#),
      565 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#06#),
      577 => to_slv(opcode_type, 16#07#),
      578 => to_slv(opcode_type, 16#05#),
      579 => to_slv(opcode_type, 16#05#),
      580 => to_slv(opcode_type, 16#11#),
      581 => to_slv(opcode_type, 16#05#),
      582 => to_slv(opcode_type, 16#04#),
      583 => to_slv(opcode_type, 16#0A#),
      584 => to_slv(opcode_type, 16#06#),
      585 => to_slv(opcode_type, 16#09#),
      586 => to_slv(opcode_type, 16#08#),
      587 => to_slv(opcode_type, 16#10#),
      588 => to_slv(opcode_type, 16#0E#),
      589 => to_slv(opcode_type, 16#07#),
      590 => to_slv(opcode_type, 16#0C#),
      591 => to_slv(opcode_type, 16#0F#),
      592 => to_slv(opcode_type, 16#07#),
      593 => to_slv(opcode_type, 16#05#),
      594 => to_slv(opcode_type, 16#0C#),
      595 => to_slv(opcode_type, 16#04#),
      596 => to_slv(opcode_type, 16#0C#),
      597 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#08#),
      609 => to_slv(opcode_type, 16#03#),
      610 => to_slv(opcode_type, 16#05#),
      611 => to_slv(opcode_type, 16#06#),
      612 => to_slv(opcode_type, 16#BD#),
      613 => to_slv(opcode_type, 16#11#),
      614 => to_slv(opcode_type, 16#06#),
      615 => to_slv(opcode_type, 16#07#),
      616 => to_slv(opcode_type, 16#09#),
      617 => to_slv(opcode_type, 16#0D#),
      618 => to_slv(opcode_type, 16#10#),
      619 => to_slv(opcode_type, 16#08#),
      620 => to_slv(opcode_type, 16#0A#),
      621 => to_slv(opcode_type, 16#0C#),
      622 => to_slv(opcode_type, 16#08#),
      623 => to_slv(opcode_type, 16#06#),
      624 => to_slv(opcode_type, 16#0D#),
      625 => to_slv(opcode_type, 16#0D#),
      626 => to_slv(opcode_type, 16#06#),
      627 => to_slv(opcode_type, 16#0D#),
      628 => to_slv(opcode_type, 16#0B#),
      629 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#08#),
      641 => to_slv(opcode_type, 16#07#),
      642 => to_slv(opcode_type, 16#02#),
      643 => to_slv(opcode_type, 16#01#),
      644 => to_slv(opcode_type, 16#0A#),
      645 => to_slv(opcode_type, 16#05#),
      646 => to_slv(opcode_type, 16#09#),
      647 => to_slv(opcode_type, 16#11#),
      648 => to_slv(opcode_type, 16#0A#),
      649 => to_slv(opcode_type, 16#09#),
      650 => to_slv(opcode_type, 16#07#),
      651 => to_slv(opcode_type, 16#05#),
      652 => to_slv(opcode_type, 16#8B#),
      653 => to_slv(opcode_type, 16#09#),
      654 => to_slv(opcode_type, 16#0E#),
      655 => to_slv(opcode_type, 16#11#),
      656 => to_slv(opcode_type, 16#06#),
      657 => to_slv(opcode_type, 16#07#),
      658 => to_slv(opcode_type, 16#11#),
      659 => to_slv(opcode_type, 16#0B#),
      660 => to_slv(opcode_type, 16#10#),
      661 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#06#),
      673 => to_slv(opcode_type, 16#06#),
      674 => to_slv(opcode_type, 16#06#),
      675 => to_slv(opcode_type, 16#06#),
      676 => to_slv(opcode_type, 16#10#),
      677 => to_slv(opcode_type, 16#0B#),
      678 => to_slv(opcode_type, 16#05#),
      679 => to_slv(opcode_type, 16#F1#),
      680 => to_slv(opcode_type, 16#01#),
      681 => to_slv(opcode_type, 16#05#),
      682 => to_slv(opcode_type, 16#18#),
      683 => to_slv(opcode_type, 16#07#),
      684 => to_slv(opcode_type, 16#02#),
      685 => to_slv(opcode_type, 16#06#),
      686 => to_slv(opcode_type, 16#0C#),
      687 => to_slv(opcode_type, 16#0C#),
      688 => to_slv(opcode_type, 16#08#),
      689 => to_slv(opcode_type, 16#09#),
      690 => to_slv(opcode_type, 16#0A#),
      691 => to_slv(opcode_type, 16#0C#),
      692 => to_slv(opcode_type, 16#0C#),
      693 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#06#),
      705 => to_slv(opcode_type, 16#09#),
      706 => to_slv(opcode_type, 16#01#),
      707 => to_slv(opcode_type, 16#02#),
      708 => to_slv(opcode_type, 16#0A#),
      709 => to_slv(opcode_type, 16#02#),
      710 => to_slv(opcode_type, 16#03#),
      711 => to_slv(opcode_type, 16#0A#),
      712 => to_slv(opcode_type, 16#07#),
      713 => to_slv(opcode_type, 16#06#),
      714 => to_slv(opcode_type, 16#02#),
      715 => to_slv(opcode_type, 16#10#),
      716 => to_slv(opcode_type, 16#02#),
      717 => to_slv(opcode_type, 16#11#),
      718 => to_slv(opcode_type, 16#07#),
      719 => to_slv(opcode_type, 16#07#),
      720 => to_slv(opcode_type, 16#0A#),
      721 => to_slv(opcode_type, 16#0D#),
      722 => to_slv(opcode_type, 16#07#),
      723 => to_slv(opcode_type, 16#0C#),
      724 => to_slv(opcode_type, 16#0F#),
      725 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#09#),
      737 => to_slv(opcode_type, 16#05#),
      738 => to_slv(opcode_type, 16#04#),
      739 => to_slv(opcode_type, 16#06#),
      740 => to_slv(opcode_type, 16#0C#),
      741 => to_slv(opcode_type, 16#0F#),
      742 => to_slv(opcode_type, 16#09#),
      743 => to_slv(opcode_type, 16#06#),
      744 => to_slv(opcode_type, 16#08#),
      745 => to_slv(opcode_type, 16#0E#),
      746 => to_slv(opcode_type, 16#0A#),
      747 => to_slv(opcode_type, 16#08#),
      748 => to_slv(opcode_type, 16#0D#),
      749 => to_slv(opcode_type, 16#11#),
      750 => to_slv(opcode_type, 16#08#),
      751 => to_slv(opcode_type, 16#08#),
      752 => to_slv(opcode_type, 16#0E#),
      753 => to_slv(opcode_type, 16#0A#),
      754 => to_slv(opcode_type, 16#09#),
      755 => to_slv(opcode_type, 16#11#),
      756 => to_slv(opcode_type, 16#10#),
      757 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#06#),
      769 => to_slv(opcode_type, 16#07#),
      770 => to_slv(opcode_type, 16#06#),
      771 => to_slv(opcode_type, 16#05#),
      772 => to_slv(opcode_type, 16#0E#),
      773 => to_slv(opcode_type, 16#05#),
      774 => to_slv(opcode_type, 16#0A#),
      775 => to_slv(opcode_type, 16#08#),
      776 => to_slv(opcode_type, 16#05#),
      777 => to_slv(opcode_type, 16#0F#),
      778 => to_slv(opcode_type, 16#01#),
      779 => to_slv(opcode_type, 16#0B#),
      780 => to_slv(opcode_type, 16#09#),
      781 => to_slv(opcode_type, 16#08#),
      782 => to_slv(opcode_type, 16#01#),
      783 => to_slv(opcode_type, 16#0E#),
      784 => to_slv(opcode_type, 16#05#),
      785 => to_slv(opcode_type, 16#C0#),
      786 => to_slv(opcode_type, 16#04#),
      787 => to_slv(opcode_type, 16#01#),
      788 => to_slv(opcode_type, 16#0C#),
      789 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#09#),
      801 => to_slv(opcode_type, 16#08#),
      802 => to_slv(opcode_type, 16#03#),
      803 => to_slv(opcode_type, 16#04#),
      804 => to_slv(opcode_type, 16#B8#),
      805 => to_slv(opcode_type, 16#09#),
      806 => to_slv(opcode_type, 16#01#),
      807 => to_slv(opcode_type, 16#0A#),
      808 => to_slv(opcode_type, 16#07#),
      809 => to_slv(opcode_type, 16#0C#),
      810 => to_slv(opcode_type, 16#0E#),
      811 => to_slv(opcode_type, 16#07#),
      812 => to_slv(opcode_type, 16#01#),
      813 => to_slv(opcode_type, 16#04#),
      814 => to_slv(opcode_type, 16#0B#),
      815 => to_slv(opcode_type, 16#06#),
      816 => to_slv(opcode_type, 16#03#),
      817 => to_slv(opcode_type, 16#11#),
      818 => to_slv(opcode_type, 16#09#),
      819 => to_slv(opcode_type, 16#10#),
      820 => to_slv(opcode_type, 16#0B#),
      821 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#06#),
      833 => to_slv(opcode_type, 16#04#),
      834 => to_slv(opcode_type, 16#03#),
      835 => to_slv(opcode_type, 16#08#),
      836 => to_slv(opcode_type, 16#0A#),
      837 => to_slv(opcode_type, 16#0A#),
      838 => to_slv(opcode_type, 16#07#),
      839 => to_slv(opcode_type, 16#06#),
      840 => to_slv(opcode_type, 16#06#),
      841 => to_slv(opcode_type, 16#11#),
      842 => to_slv(opcode_type, 16#0C#),
      843 => to_slv(opcode_type, 16#09#),
      844 => to_slv(opcode_type, 16#10#),
      845 => to_slv(opcode_type, 16#D4#),
      846 => to_slv(opcode_type, 16#07#),
      847 => to_slv(opcode_type, 16#08#),
      848 => to_slv(opcode_type, 16#0D#),
      849 => to_slv(opcode_type, 16#11#),
      850 => to_slv(opcode_type, 16#07#),
      851 => to_slv(opcode_type, 16#11#),
      852 => to_slv(opcode_type, 16#11#),
      853 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#09#),
      865 => to_slv(opcode_type, 16#04#),
      866 => to_slv(opcode_type, 16#06#),
      867 => to_slv(opcode_type, 16#06#),
      868 => to_slv(opcode_type, 16#10#),
      869 => to_slv(opcode_type, 16#0D#),
      870 => to_slv(opcode_type, 16#03#),
      871 => to_slv(opcode_type, 16#0E#),
      872 => to_slv(opcode_type, 16#09#),
      873 => to_slv(opcode_type, 16#06#),
      874 => to_slv(opcode_type, 16#05#),
      875 => to_slv(opcode_type, 16#0C#),
      876 => to_slv(opcode_type, 16#02#),
      877 => to_slv(opcode_type, 16#0D#),
      878 => to_slv(opcode_type, 16#09#),
      879 => to_slv(opcode_type, 16#06#),
      880 => to_slv(opcode_type, 16#11#),
      881 => to_slv(opcode_type, 16#0E#),
      882 => to_slv(opcode_type, 16#08#),
      883 => to_slv(opcode_type, 16#0E#),
      884 => to_slv(opcode_type, 16#11#),
      885 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#09#),
      897 => to_slv(opcode_type, 16#09#),
      898 => to_slv(opcode_type, 16#04#),
      899 => to_slv(opcode_type, 16#01#),
      900 => to_slv(opcode_type, 16#0B#),
      901 => to_slv(opcode_type, 16#07#),
      902 => to_slv(opcode_type, 16#01#),
      903 => to_slv(opcode_type, 16#10#),
      904 => to_slv(opcode_type, 16#03#),
      905 => to_slv(opcode_type, 16#0E#),
      906 => to_slv(opcode_type, 16#07#),
      907 => to_slv(opcode_type, 16#08#),
      908 => to_slv(opcode_type, 16#07#),
      909 => to_slv(opcode_type, 16#0D#),
      910 => to_slv(opcode_type, 16#0E#),
      911 => to_slv(opcode_type, 16#07#),
      912 => to_slv(opcode_type, 16#11#),
      913 => to_slv(opcode_type, 16#0A#),
      914 => to_slv(opcode_type, 16#05#),
      915 => to_slv(opcode_type, 16#02#),
      916 => to_slv(opcode_type, 16#10#),
      917 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#09#),
      929 => to_slv(opcode_type, 16#08#),
      930 => to_slv(opcode_type, 16#06#),
      931 => to_slv(opcode_type, 16#04#),
      932 => to_slv(opcode_type, 16#0A#),
      933 => to_slv(opcode_type, 16#05#),
      934 => to_slv(opcode_type, 16#8F#),
      935 => to_slv(opcode_type, 16#09#),
      936 => to_slv(opcode_type, 16#08#),
      937 => to_slv(opcode_type, 16#0A#),
      938 => to_slv(opcode_type, 16#D6#),
      939 => to_slv(opcode_type, 16#01#),
      940 => to_slv(opcode_type, 16#0B#),
      941 => to_slv(opcode_type, 16#01#),
      942 => to_slv(opcode_type, 16#07#),
      943 => to_slv(opcode_type, 16#07#),
      944 => to_slv(opcode_type, 16#0D#),
      945 => to_slv(opcode_type, 16#0E#),
      946 => to_slv(opcode_type, 16#09#),
      947 => to_slv(opcode_type, 16#0F#),
      948 => to_slv(opcode_type, 16#0D#),
      949 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#05#),
      962 => to_slv(opcode_type, 16#03#),
      963 => to_slv(opcode_type, 16#08#),
      964 => to_slv(opcode_type, 16#0E#),
      965 => to_slv(opcode_type, 16#0E#),
      966 => to_slv(opcode_type, 16#09#),
      967 => to_slv(opcode_type, 16#09#),
      968 => to_slv(opcode_type, 16#07#),
      969 => to_slv(opcode_type, 16#0A#),
      970 => to_slv(opcode_type, 16#0B#),
      971 => to_slv(opcode_type, 16#06#),
      972 => to_slv(opcode_type, 16#0C#),
      973 => to_slv(opcode_type, 16#0F#),
      974 => to_slv(opcode_type, 16#06#),
      975 => to_slv(opcode_type, 16#07#),
      976 => to_slv(opcode_type, 16#11#),
      977 => to_slv(opcode_type, 16#10#),
      978 => to_slv(opcode_type, 16#09#),
      979 => to_slv(opcode_type, 16#0A#),
      980 => to_slv(opcode_type, 16#0C#),
      981 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#08#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#03#),
      995 => to_slv(opcode_type, 16#01#),
      996 => to_slv(opcode_type, 16#0B#),
      997 => to_slv(opcode_type, 16#04#),
      998 => to_slv(opcode_type, 16#02#),
      999 => to_slv(opcode_type, 16#48#),
      1000 => to_slv(opcode_type, 16#09#),
      1001 => to_slv(opcode_type, 16#08#),
      1002 => to_slv(opcode_type, 16#03#),
      1003 => to_slv(opcode_type, 16#0E#),
      1004 => to_slv(opcode_type, 16#09#),
      1005 => to_slv(opcode_type, 16#8B#),
      1006 => to_slv(opcode_type, 16#0F#),
      1007 => to_slv(opcode_type, 16#09#),
      1008 => to_slv(opcode_type, 16#01#),
      1009 => to_slv(opcode_type, 16#0E#),
      1010 => to_slv(opcode_type, 16#07#),
      1011 => to_slv(opcode_type, 16#CC#),
      1012 => to_slv(opcode_type, 16#0F#),
      1013 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#08#),
      1025 => to_slv(opcode_type, 16#02#),
      1026 => to_slv(opcode_type, 16#07#),
      1027 => to_slv(opcode_type, 16#05#),
      1028 => to_slv(opcode_type, 16#0E#),
      1029 => to_slv(opcode_type, 16#02#),
      1030 => to_slv(opcode_type, 16#11#),
      1031 => to_slv(opcode_type, 16#06#),
      1032 => to_slv(opcode_type, 16#08#),
      1033 => to_slv(opcode_type, 16#04#),
      1034 => to_slv(opcode_type, 16#0A#),
      1035 => to_slv(opcode_type, 16#06#),
      1036 => to_slv(opcode_type, 16#11#),
      1037 => to_slv(opcode_type, 16#10#),
      1038 => to_slv(opcode_type, 16#09#),
      1039 => to_slv(opcode_type, 16#08#),
      1040 => to_slv(opcode_type, 16#0F#),
      1041 => to_slv(opcode_type, 16#0A#),
      1042 => to_slv(opcode_type, 16#09#),
      1043 => to_slv(opcode_type, 16#6E#),
      1044 => to_slv(opcode_type, 16#0B#),
      1045 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#08#),
      1057 => to_slv(opcode_type, 16#01#),
      1058 => to_slv(opcode_type, 16#09#),
      1059 => to_slv(opcode_type, 16#06#),
      1060 => to_slv(opcode_type, 16#32#),
      1061 => to_slv(opcode_type, 16#0E#),
      1062 => to_slv(opcode_type, 16#09#),
      1063 => to_slv(opcode_type, 16#0B#),
      1064 => to_slv(opcode_type, 16#10#),
      1065 => to_slv(opcode_type, 16#07#),
      1066 => to_slv(opcode_type, 16#02#),
      1067 => to_slv(opcode_type, 16#06#),
      1068 => to_slv(opcode_type, 16#0D#),
      1069 => to_slv(opcode_type, 16#0F#),
      1070 => to_slv(opcode_type, 16#09#),
      1071 => to_slv(opcode_type, 16#08#),
      1072 => to_slv(opcode_type, 16#0E#),
      1073 => to_slv(opcode_type, 16#E5#),
      1074 => to_slv(opcode_type, 16#07#),
      1075 => to_slv(opcode_type, 16#E3#),
      1076 => to_slv(opcode_type, 16#0B#),
      1077 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#08#),
      1089 => to_slv(opcode_type, 16#04#),
      1090 => to_slv(opcode_type, 16#09#),
      1091 => to_slv(opcode_type, 16#01#),
      1092 => to_slv(opcode_type, 16#10#),
      1093 => to_slv(opcode_type, 16#05#),
      1094 => to_slv(opcode_type, 16#0B#),
      1095 => to_slv(opcode_type, 16#09#),
      1096 => to_slv(opcode_type, 16#09#),
      1097 => to_slv(opcode_type, 16#07#),
      1098 => to_slv(opcode_type, 16#0F#),
      1099 => to_slv(opcode_type, 16#0B#),
      1100 => to_slv(opcode_type, 16#09#),
      1101 => to_slv(opcode_type, 16#0E#),
      1102 => to_slv(opcode_type, 16#0F#),
      1103 => to_slv(opcode_type, 16#09#),
      1104 => to_slv(opcode_type, 16#07#),
      1105 => to_slv(opcode_type, 16#12#),
      1106 => to_slv(opcode_type, 16#27#),
      1107 => to_slv(opcode_type, 16#03#),
      1108 => to_slv(opcode_type, 16#0D#),
      1109 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#07#),
      1121 => to_slv(opcode_type, 16#03#),
      1122 => to_slv(opcode_type, 16#06#),
      1123 => to_slv(opcode_type, 16#04#),
      1124 => to_slv(opcode_type, 16#11#),
      1125 => to_slv(opcode_type, 16#08#),
      1126 => to_slv(opcode_type, 16#0D#),
      1127 => to_slv(opcode_type, 16#0B#),
      1128 => to_slv(opcode_type, 16#09#),
      1129 => to_slv(opcode_type, 16#07#),
      1130 => to_slv(opcode_type, 16#01#),
      1131 => to_slv(opcode_type, 16#0D#),
      1132 => to_slv(opcode_type, 16#03#),
      1133 => to_slv(opcode_type, 16#11#),
      1134 => to_slv(opcode_type, 16#09#),
      1135 => to_slv(opcode_type, 16#08#),
      1136 => to_slv(opcode_type, 16#0A#),
      1137 => to_slv(opcode_type, 16#0D#),
      1138 => to_slv(opcode_type, 16#07#),
      1139 => to_slv(opcode_type, 16#10#),
      1140 => to_slv(opcode_type, 16#0C#),
      1141 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#08#),
      1153 => to_slv(opcode_type, 16#01#),
      1154 => to_slv(opcode_type, 16#09#),
      1155 => to_slv(opcode_type, 16#07#),
      1156 => to_slv(opcode_type, 16#0F#),
      1157 => to_slv(opcode_type, 16#10#),
      1158 => to_slv(opcode_type, 16#05#),
      1159 => to_slv(opcode_type, 16#11#),
      1160 => to_slv(opcode_type, 16#06#),
      1161 => to_slv(opcode_type, 16#06#),
      1162 => to_slv(opcode_type, 16#04#),
      1163 => to_slv(opcode_type, 16#0E#),
      1164 => to_slv(opcode_type, 16#03#),
      1165 => to_slv(opcode_type, 16#0B#),
      1166 => to_slv(opcode_type, 16#08#),
      1167 => to_slv(opcode_type, 16#07#),
      1168 => to_slv(opcode_type, 16#0A#),
      1169 => to_slv(opcode_type, 16#10#),
      1170 => to_slv(opcode_type, 16#09#),
      1171 => to_slv(opcode_type, 16#0E#),
      1172 => to_slv(opcode_type, 16#81#),
      1173 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#08#),
      1185 => to_slv(opcode_type, 16#06#),
      1186 => to_slv(opcode_type, 16#05#),
      1187 => to_slv(opcode_type, 16#03#),
      1188 => to_slv(opcode_type, 16#0C#),
      1189 => to_slv(opcode_type, 16#05#),
      1190 => to_slv(opcode_type, 16#01#),
      1191 => to_slv(opcode_type, 16#C7#),
      1192 => to_slv(opcode_type, 16#09#),
      1193 => to_slv(opcode_type, 16#08#),
      1194 => to_slv(opcode_type, 16#04#),
      1195 => to_slv(opcode_type, 16#3A#),
      1196 => to_slv(opcode_type, 16#02#),
      1197 => to_slv(opcode_type, 16#10#),
      1198 => to_slv(opcode_type, 16#07#),
      1199 => to_slv(opcode_type, 16#09#),
      1200 => to_slv(opcode_type, 16#0B#),
      1201 => to_slv(opcode_type, 16#10#),
      1202 => to_slv(opcode_type, 16#06#),
      1203 => to_slv(opcode_type, 16#0B#),
      1204 => to_slv(opcode_type, 16#0D#),
      1205 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#07#),
      1217 => to_slv(opcode_type, 16#03#),
      1218 => to_slv(opcode_type, 16#05#),
      1219 => to_slv(opcode_type, 16#09#),
      1220 => to_slv(opcode_type, 16#0D#),
      1221 => to_slv(opcode_type, 16#0B#),
      1222 => to_slv(opcode_type, 16#09#),
      1223 => to_slv(opcode_type, 16#09#),
      1224 => to_slv(opcode_type, 16#08#),
      1225 => to_slv(opcode_type, 16#7C#),
      1226 => to_slv(opcode_type, 16#0F#),
      1227 => to_slv(opcode_type, 16#07#),
      1228 => to_slv(opcode_type, 16#0B#),
      1229 => to_slv(opcode_type, 16#0C#),
      1230 => to_slv(opcode_type, 16#08#),
      1231 => to_slv(opcode_type, 16#06#),
      1232 => to_slv(opcode_type, 16#0A#),
      1233 => to_slv(opcode_type, 16#0F#),
      1234 => to_slv(opcode_type, 16#08#),
      1235 => to_slv(opcode_type, 16#0D#),
      1236 => to_slv(opcode_type, 16#0D#),
      1237 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#06#),
      1249 => to_slv(opcode_type, 16#08#),
      1250 => to_slv(opcode_type, 16#03#),
      1251 => to_slv(opcode_type, 16#01#),
      1252 => to_slv(opcode_type, 16#0E#),
      1253 => to_slv(opcode_type, 16#05#),
      1254 => to_slv(opcode_type, 16#02#),
      1255 => to_slv(opcode_type, 16#10#),
      1256 => to_slv(opcode_type, 16#08#),
      1257 => to_slv(opcode_type, 16#07#),
      1258 => to_slv(opcode_type, 16#02#),
      1259 => to_slv(opcode_type, 16#0E#),
      1260 => to_slv(opcode_type, 16#06#),
      1261 => to_slv(opcode_type, 16#0A#),
      1262 => to_slv(opcode_type, 16#0B#),
      1263 => to_slv(opcode_type, 16#09#),
      1264 => to_slv(opcode_type, 16#04#),
      1265 => to_slv(opcode_type, 16#0D#),
      1266 => to_slv(opcode_type, 16#07#),
      1267 => to_slv(opcode_type, 16#10#),
      1268 => to_slv(opcode_type, 16#0A#),
      1269 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#01#),
      1282 => to_slv(opcode_type, 16#08#),
      1283 => to_slv(opcode_type, 16#06#),
      1284 => to_slv(opcode_type, 16#75#),
      1285 => to_slv(opcode_type, 16#0D#),
      1286 => to_slv(opcode_type, 16#07#),
      1287 => to_slv(opcode_type, 16#0E#),
      1288 => to_slv(opcode_type, 16#0E#),
      1289 => to_slv(opcode_type, 16#06#),
      1290 => to_slv(opcode_type, 16#03#),
      1291 => to_slv(opcode_type, 16#06#),
      1292 => to_slv(opcode_type, 16#0E#),
      1293 => to_slv(opcode_type, 16#0D#),
      1294 => to_slv(opcode_type, 16#09#),
      1295 => to_slv(opcode_type, 16#07#),
      1296 => to_slv(opcode_type, 16#0F#),
      1297 => to_slv(opcode_type, 16#87#),
      1298 => to_slv(opcode_type, 16#08#),
      1299 => to_slv(opcode_type, 16#10#),
      1300 => to_slv(opcode_type, 16#0D#),
      1301 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#08#),
      1313 => to_slv(opcode_type, 16#03#),
      1314 => to_slv(opcode_type, 16#09#),
      1315 => to_slv(opcode_type, 16#07#),
      1316 => to_slv(opcode_type, 16#0F#),
      1317 => to_slv(opcode_type, 16#0D#),
      1318 => to_slv(opcode_type, 16#01#),
      1319 => to_slv(opcode_type, 16#0D#),
      1320 => to_slv(opcode_type, 16#09#),
      1321 => to_slv(opcode_type, 16#06#),
      1322 => to_slv(opcode_type, 16#09#),
      1323 => to_slv(opcode_type, 16#10#),
      1324 => to_slv(opcode_type, 16#0E#),
      1325 => to_slv(opcode_type, 16#08#),
      1326 => to_slv(opcode_type, 16#0B#),
      1327 => to_slv(opcode_type, 16#11#),
      1328 => to_slv(opcode_type, 16#08#),
      1329 => to_slv(opcode_type, 16#03#),
      1330 => to_slv(opcode_type, 16#0F#),
      1331 => to_slv(opcode_type, 16#04#),
      1332 => to_slv(opcode_type, 16#0C#),
      1333 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#08#),
      1345 => to_slv(opcode_type, 16#04#),
      1346 => to_slv(opcode_type, 16#05#),
      1347 => to_slv(opcode_type, 16#06#),
      1348 => to_slv(opcode_type, 16#11#),
      1349 => to_slv(opcode_type, 16#11#),
      1350 => to_slv(opcode_type, 16#09#),
      1351 => to_slv(opcode_type, 16#07#),
      1352 => to_slv(opcode_type, 16#07#),
      1353 => to_slv(opcode_type, 16#11#),
      1354 => to_slv(opcode_type, 16#F4#),
      1355 => to_slv(opcode_type, 16#08#),
      1356 => to_slv(opcode_type, 16#0D#),
      1357 => to_slv(opcode_type, 16#0D#),
      1358 => to_slv(opcode_type, 16#06#),
      1359 => to_slv(opcode_type, 16#07#),
      1360 => to_slv(opcode_type, 16#B9#),
      1361 => to_slv(opcode_type, 16#0B#),
      1362 => to_slv(opcode_type, 16#07#),
      1363 => to_slv(opcode_type, 16#0E#),
      1364 => to_slv(opcode_type, 16#11#),
      1365 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#06#),
      1377 => to_slv(opcode_type, 16#09#),
      1378 => to_slv(opcode_type, 16#03#),
      1379 => to_slv(opcode_type, 16#09#),
      1380 => to_slv(opcode_type, 16#9D#),
      1381 => to_slv(opcode_type, 16#0F#),
      1382 => to_slv(opcode_type, 16#01#),
      1383 => to_slv(opcode_type, 16#01#),
      1384 => to_slv(opcode_type, 16#0A#),
      1385 => to_slv(opcode_type, 16#09#),
      1386 => to_slv(opcode_type, 16#04#),
      1387 => to_slv(opcode_type, 16#07#),
      1388 => to_slv(opcode_type, 16#0E#),
      1389 => to_slv(opcode_type, 16#10#),
      1390 => to_slv(opcode_type, 16#08#),
      1391 => to_slv(opcode_type, 16#08#),
      1392 => to_slv(opcode_type, 16#10#),
      1393 => to_slv(opcode_type, 16#0C#),
      1394 => to_slv(opcode_type, 16#09#),
      1395 => to_slv(opcode_type, 16#0E#),
      1396 => to_slv(opcode_type, 16#0B#),
      1397 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#09#),
      1409 => to_slv(opcode_type, 16#08#),
      1410 => to_slv(opcode_type, 16#09#),
      1411 => to_slv(opcode_type, 16#09#),
      1412 => to_slv(opcode_type, 16#11#),
      1413 => to_slv(opcode_type, 16#10#),
      1414 => to_slv(opcode_type, 16#06#),
      1415 => to_slv(opcode_type, 16#0F#),
      1416 => to_slv(opcode_type, 16#0E#),
      1417 => to_slv(opcode_type, 16#01#),
      1418 => to_slv(opcode_type, 16#06#),
      1419 => to_slv(opcode_type, 16#0C#),
      1420 => to_slv(opcode_type, 16#0A#),
      1421 => to_slv(opcode_type, 16#04#),
      1422 => to_slv(opcode_type, 16#09#),
      1423 => to_slv(opcode_type, 16#08#),
      1424 => to_slv(opcode_type, 16#0E#),
      1425 => to_slv(opcode_type, 16#0D#),
      1426 => to_slv(opcode_type, 16#07#),
      1427 => to_slv(opcode_type, 16#0E#),
      1428 => to_slv(opcode_type, 16#0C#),
      1429 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#07#),
      1441 => to_slv(opcode_type, 16#04#),
      1442 => to_slv(opcode_type, 16#09#),
      1443 => to_slv(opcode_type, 16#07#),
      1444 => to_slv(opcode_type, 16#0D#),
      1445 => to_slv(opcode_type, 16#0B#),
      1446 => to_slv(opcode_type, 16#04#),
      1447 => to_slv(opcode_type, 16#0D#),
      1448 => to_slv(opcode_type, 16#06#),
      1449 => to_slv(opcode_type, 16#07#),
      1450 => to_slv(opcode_type, 16#09#),
      1451 => to_slv(opcode_type, 16#0A#),
      1452 => to_slv(opcode_type, 16#0F#),
      1453 => to_slv(opcode_type, 16#06#),
      1454 => to_slv(opcode_type, 16#0A#),
      1455 => to_slv(opcode_type, 16#11#),
      1456 => to_slv(opcode_type, 16#09#),
      1457 => to_slv(opcode_type, 16#08#),
      1458 => to_slv(opcode_type, 16#0B#),
      1459 => to_slv(opcode_type, 16#0C#),
      1460 => to_slv(opcode_type, 16#11#),
      1461 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#07#),
      1473 => to_slv(opcode_type, 16#04#),
      1474 => to_slv(opcode_type, 16#01#),
      1475 => to_slv(opcode_type, 16#06#),
      1476 => to_slv(opcode_type, 16#67#),
      1477 => to_slv(opcode_type, 16#0C#),
      1478 => to_slv(opcode_type, 16#07#),
      1479 => to_slv(opcode_type, 16#09#),
      1480 => to_slv(opcode_type, 16#07#),
      1481 => to_slv(opcode_type, 16#0C#),
      1482 => to_slv(opcode_type, 16#0A#),
      1483 => to_slv(opcode_type, 16#08#),
      1484 => to_slv(opcode_type, 16#11#),
      1485 => to_slv(opcode_type, 16#0F#),
      1486 => to_slv(opcode_type, 16#08#),
      1487 => to_slv(opcode_type, 16#06#),
      1488 => to_slv(opcode_type, 16#0A#),
      1489 => to_slv(opcode_type, 16#0E#),
      1490 => to_slv(opcode_type, 16#06#),
      1491 => to_slv(opcode_type, 16#0F#),
      1492 => to_slv(opcode_type, 16#11#),
      1493 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#06#),
      1505 => to_slv(opcode_type, 16#04#),
      1506 => to_slv(opcode_type, 16#02#),
      1507 => to_slv(opcode_type, 16#07#),
      1508 => to_slv(opcode_type, 16#DE#),
      1509 => to_slv(opcode_type, 16#0C#),
      1510 => to_slv(opcode_type, 16#09#),
      1511 => to_slv(opcode_type, 16#07#),
      1512 => to_slv(opcode_type, 16#08#),
      1513 => to_slv(opcode_type, 16#0A#),
      1514 => to_slv(opcode_type, 16#0A#),
      1515 => to_slv(opcode_type, 16#08#),
      1516 => to_slv(opcode_type, 16#0E#),
      1517 => to_slv(opcode_type, 16#0A#),
      1518 => to_slv(opcode_type, 16#09#),
      1519 => to_slv(opcode_type, 16#09#),
      1520 => to_slv(opcode_type, 16#0D#),
      1521 => to_slv(opcode_type, 16#0C#),
      1522 => to_slv(opcode_type, 16#07#),
      1523 => to_slv(opcode_type, 16#10#),
      1524 => to_slv(opcode_type, 16#DC#),
      1525 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#09#),
      1537 => to_slv(opcode_type, 16#01#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#08#),
      1540 => to_slv(opcode_type, 16#0D#),
      1541 => to_slv(opcode_type, 16#0A#),
      1542 => to_slv(opcode_type, 16#09#),
      1543 => to_slv(opcode_type, 16#10#),
      1544 => to_slv(opcode_type, 16#0B#),
      1545 => to_slv(opcode_type, 16#07#),
      1546 => to_slv(opcode_type, 16#04#),
      1547 => to_slv(opcode_type, 16#09#),
      1548 => to_slv(opcode_type, 16#0B#),
      1549 => to_slv(opcode_type, 16#0F#),
      1550 => to_slv(opcode_type, 16#06#),
      1551 => to_slv(opcode_type, 16#09#),
      1552 => to_slv(opcode_type, 16#0A#),
      1553 => to_slv(opcode_type, 16#0F#),
      1554 => to_slv(opcode_type, 16#09#),
      1555 => to_slv(opcode_type, 16#0B#),
      1556 => to_slv(opcode_type, 16#0A#),
      1557 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#09#),
      1569 => to_slv(opcode_type, 16#06#),
      1570 => to_slv(opcode_type, 16#05#),
      1571 => to_slv(opcode_type, 16#06#),
      1572 => to_slv(opcode_type, 16#0F#),
      1573 => to_slv(opcode_type, 16#0C#),
      1574 => to_slv(opcode_type, 16#01#),
      1575 => to_slv(opcode_type, 16#02#),
      1576 => to_slv(opcode_type, 16#0D#),
      1577 => to_slv(opcode_type, 16#07#),
      1578 => to_slv(opcode_type, 16#08#),
      1579 => to_slv(opcode_type, 16#01#),
      1580 => to_slv(opcode_type, 16#0B#),
      1581 => to_slv(opcode_type, 16#02#),
      1582 => to_slv(opcode_type, 16#0D#),
      1583 => to_slv(opcode_type, 16#06#),
      1584 => to_slv(opcode_type, 16#08#),
      1585 => to_slv(opcode_type, 16#0A#),
      1586 => to_slv(opcode_type, 16#10#),
      1587 => to_slv(opcode_type, 16#02#),
      1588 => to_slv(opcode_type, 16#0E#),
      1589 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#07#),
      1601 => to_slv(opcode_type, 16#02#),
      1602 => to_slv(opcode_type, 16#07#),
      1603 => to_slv(opcode_type, 16#02#),
      1604 => to_slv(opcode_type, 16#76#),
      1605 => to_slv(opcode_type, 16#08#),
      1606 => to_slv(opcode_type, 16#0F#),
      1607 => to_slv(opcode_type, 16#11#),
      1608 => to_slv(opcode_type, 16#07#),
      1609 => to_slv(opcode_type, 16#09#),
      1610 => to_slv(opcode_type, 16#01#),
      1611 => to_slv(opcode_type, 16#0F#),
      1612 => to_slv(opcode_type, 16#05#),
      1613 => to_slv(opcode_type, 16#CB#),
      1614 => to_slv(opcode_type, 16#06#),
      1615 => to_slv(opcode_type, 16#06#),
      1616 => to_slv(opcode_type, 16#93#),
      1617 => to_slv(opcode_type, 16#0E#),
      1618 => to_slv(opcode_type, 16#06#),
      1619 => to_slv(opcode_type, 16#0B#),
      1620 => to_slv(opcode_type, 16#0E#),
      1621 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#07#),
      1633 => to_slv(opcode_type, 16#08#),
      1634 => to_slv(opcode_type, 16#06#),
      1635 => to_slv(opcode_type, 16#04#),
      1636 => to_slv(opcode_type, 16#9B#),
      1637 => to_slv(opcode_type, 16#01#),
      1638 => to_slv(opcode_type, 16#10#),
      1639 => to_slv(opcode_type, 16#04#),
      1640 => to_slv(opcode_type, 16#07#),
      1641 => to_slv(opcode_type, 16#0E#),
      1642 => to_slv(opcode_type, 16#0E#),
      1643 => to_slv(opcode_type, 16#06#),
      1644 => to_slv(opcode_type, 16#05#),
      1645 => to_slv(opcode_type, 16#03#),
      1646 => to_slv(opcode_type, 16#10#),
      1647 => to_slv(opcode_type, 16#06#),
      1648 => to_slv(opcode_type, 16#03#),
      1649 => to_slv(opcode_type, 16#DC#),
      1650 => to_slv(opcode_type, 16#06#),
      1651 => to_slv(opcode_type, 16#0C#),
      1652 => to_slv(opcode_type, 16#0B#),
      1653 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#06#),
      1665 => to_slv(opcode_type, 16#06#),
      1666 => to_slv(opcode_type, 16#06#),
      1667 => to_slv(opcode_type, 16#01#),
      1668 => to_slv(opcode_type, 16#0E#),
      1669 => to_slv(opcode_type, 16#08#),
      1670 => to_slv(opcode_type, 16#CB#),
      1671 => to_slv(opcode_type, 16#10#),
      1672 => to_slv(opcode_type, 16#08#),
      1673 => to_slv(opcode_type, 16#09#),
      1674 => to_slv(opcode_type, 16#9C#),
      1675 => to_slv(opcode_type, 16#0F#),
      1676 => to_slv(opcode_type, 16#08#),
      1677 => to_slv(opcode_type, 16#0C#),
      1678 => to_slv(opcode_type, 16#0D#),
      1679 => to_slv(opcode_type, 16#07#),
      1680 => to_slv(opcode_type, 16#08#),
      1681 => to_slv(opcode_type, 16#05#),
      1682 => to_slv(opcode_type, 16#0F#),
      1683 => to_slv(opcode_type, 16#0B#),
      1684 => to_slv(opcode_type, 16#0C#),
      1685 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#07#),
      1697 => to_slv(opcode_type, 16#06#),
      1698 => to_slv(opcode_type, 16#01#),
      1699 => to_slv(opcode_type, 16#03#),
      1700 => to_slv(opcode_type, 16#0F#),
      1701 => to_slv(opcode_type, 16#01#),
      1702 => to_slv(opcode_type, 16#01#),
      1703 => to_slv(opcode_type, 16#11#),
      1704 => to_slv(opcode_type, 16#08#),
      1705 => to_slv(opcode_type, 16#07#),
      1706 => to_slv(opcode_type, 16#08#),
      1707 => to_slv(opcode_type, 16#11#),
      1708 => to_slv(opcode_type, 16#0A#),
      1709 => to_slv(opcode_type, 16#04#),
      1710 => to_slv(opcode_type, 16#0D#),
      1711 => to_slv(opcode_type, 16#07#),
      1712 => to_slv(opcode_type, 16#07#),
      1713 => to_slv(opcode_type, 16#0A#),
      1714 => to_slv(opcode_type, 16#0F#),
      1715 => to_slv(opcode_type, 16#03#),
      1716 => to_slv(opcode_type, 16#0A#),
      1717 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#06#),
      1729 => to_slv(opcode_type, 16#01#),
      1730 => to_slv(opcode_type, 16#06#),
      1731 => to_slv(opcode_type, 16#04#),
      1732 => to_slv(opcode_type, 16#0A#),
      1733 => to_slv(opcode_type, 16#07#),
      1734 => to_slv(opcode_type, 16#0E#),
      1735 => to_slv(opcode_type, 16#0A#),
      1736 => to_slv(opcode_type, 16#06#),
      1737 => to_slv(opcode_type, 16#06#),
      1738 => to_slv(opcode_type, 16#07#),
      1739 => to_slv(opcode_type, 16#0B#),
      1740 => to_slv(opcode_type, 16#10#),
      1741 => to_slv(opcode_type, 16#01#),
      1742 => to_slv(opcode_type, 16#11#),
      1743 => to_slv(opcode_type, 16#09#),
      1744 => to_slv(opcode_type, 16#03#),
      1745 => to_slv(opcode_type, 16#0C#),
      1746 => to_slv(opcode_type, 16#06#),
      1747 => to_slv(opcode_type, 16#B2#),
      1748 => to_slv(opcode_type, 16#40#),
      1749 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#08#),
      1761 => to_slv(opcode_type, 16#03#),
      1762 => to_slv(opcode_type, 16#02#),
      1763 => to_slv(opcode_type, 16#07#),
      1764 => to_slv(opcode_type, 16#10#),
      1765 => to_slv(opcode_type, 16#0A#),
      1766 => to_slv(opcode_type, 16#08#),
      1767 => to_slv(opcode_type, 16#09#),
      1768 => to_slv(opcode_type, 16#08#),
      1769 => to_slv(opcode_type, 16#0E#),
      1770 => to_slv(opcode_type, 16#10#),
      1771 => to_slv(opcode_type, 16#09#),
      1772 => to_slv(opcode_type, 16#0B#),
      1773 => to_slv(opcode_type, 16#0E#),
      1774 => to_slv(opcode_type, 16#09#),
      1775 => to_slv(opcode_type, 16#08#),
      1776 => to_slv(opcode_type, 16#0C#),
      1777 => to_slv(opcode_type, 16#0A#),
      1778 => to_slv(opcode_type, 16#07#),
      1779 => to_slv(opcode_type, 16#0F#),
      1780 => to_slv(opcode_type, 16#0D#),
      1781 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#07#),
      1793 => to_slv(opcode_type, 16#06#),
      1794 => to_slv(opcode_type, 16#09#),
      1795 => to_slv(opcode_type, 16#06#),
      1796 => to_slv(opcode_type, 16#0C#),
      1797 => to_slv(opcode_type, 16#11#),
      1798 => to_slv(opcode_type, 16#07#),
      1799 => to_slv(opcode_type, 16#0D#),
      1800 => to_slv(opcode_type, 16#11#),
      1801 => to_slv(opcode_type, 16#09#),
      1802 => to_slv(opcode_type, 16#08#),
      1803 => to_slv(opcode_type, 16#0E#),
      1804 => to_slv(opcode_type, 16#0B#),
      1805 => to_slv(opcode_type, 16#04#),
      1806 => to_slv(opcode_type, 16#10#),
      1807 => to_slv(opcode_type, 16#01#),
      1808 => to_slv(opcode_type, 16#06#),
      1809 => to_slv(opcode_type, 16#02#),
      1810 => to_slv(opcode_type, 16#0E#),
      1811 => to_slv(opcode_type, 16#03#),
      1812 => to_slv(opcode_type, 16#0A#),
      1813 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#08#),
      1825 => to_slv(opcode_type, 16#01#),
      1826 => to_slv(opcode_type, 16#09#),
      1827 => to_slv(opcode_type, 16#09#),
      1828 => to_slv(opcode_type, 16#0C#),
      1829 => to_slv(opcode_type, 16#11#),
      1830 => to_slv(opcode_type, 16#06#),
      1831 => to_slv(opcode_type, 16#A2#),
      1832 => to_slv(opcode_type, 16#0A#),
      1833 => to_slv(opcode_type, 16#08#),
      1834 => to_slv(opcode_type, 16#03#),
      1835 => to_slv(opcode_type, 16#08#),
      1836 => to_slv(opcode_type, 16#11#),
      1837 => to_slv(opcode_type, 16#AF#),
      1838 => to_slv(opcode_type, 16#08#),
      1839 => to_slv(opcode_type, 16#08#),
      1840 => to_slv(opcode_type, 16#0F#),
      1841 => to_slv(opcode_type, 16#10#),
      1842 => to_slv(opcode_type, 16#08#),
      1843 => to_slv(opcode_type, 16#10#),
      1844 => to_slv(opcode_type, 16#0B#),
      1845 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#06#),
      1857 => to_slv(opcode_type, 16#06#),
      1858 => to_slv(opcode_type, 16#07#),
      1859 => to_slv(opcode_type, 16#05#),
      1860 => to_slv(opcode_type, 16#0D#),
      1861 => to_slv(opcode_type, 16#03#),
      1862 => to_slv(opcode_type, 16#0F#),
      1863 => to_slv(opcode_type, 16#06#),
      1864 => to_slv(opcode_type, 16#09#),
      1865 => to_slv(opcode_type, 16#0E#),
      1866 => to_slv(opcode_type, 16#0F#),
      1867 => to_slv(opcode_type, 16#01#),
      1868 => to_slv(opcode_type, 16#11#),
      1869 => to_slv(opcode_type, 16#04#),
      1870 => to_slv(opcode_type, 16#07#),
      1871 => to_slv(opcode_type, 16#07#),
      1872 => to_slv(opcode_type, 16#0E#),
      1873 => to_slv(opcode_type, 16#10#),
      1874 => to_slv(opcode_type, 16#07#),
      1875 => to_slv(opcode_type, 16#0D#),
      1876 => to_slv(opcode_type, 16#96#),
      1877 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#08#),
      1889 => to_slv(opcode_type, 16#02#),
      1890 => to_slv(opcode_type, 16#07#),
      1891 => to_slv(opcode_type, 16#08#),
      1892 => to_slv(opcode_type, 16#59#),
      1893 => to_slv(opcode_type, 16#10#),
      1894 => to_slv(opcode_type, 16#01#),
      1895 => to_slv(opcode_type, 16#0B#),
      1896 => to_slv(opcode_type, 16#08#),
      1897 => to_slv(opcode_type, 16#08#),
      1898 => to_slv(opcode_type, 16#03#),
      1899 => to_slv(opcode_type, 16#80#),
      1900 => to_slv(opcode_type, 16#01#),
      1901 => to_slv(opcode_type, 16#3F#),
      1902 => to_slv(opcode_type, 16#07#),
      1903 => to_slv(opcode_type, 16#07#),
      1904 => to_slv(opcode_type, 16#11#),
      1905 => to_slv(opcode_type, 16#10#),
      1906 => to_slv(opcode_type, 16#06#),
      1907 => to_slv(opcode_type, 16#0A#),
      1908 => to_slv(opcode_type, 16#11#),
      1909 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#07#),
      1921 => to_slv(opcode_type, 16#05#),
      1922 => to_slv(opcode_type, 16#01#),
      1923 => to_slv(opcode_type, 16#09#),
      1924 => to_slv(opcode_type, 16#0F#),
      1925 => to_slv(opcode_type, 16#0F#),
      1926 => to_slv(opcode_type, 16#09#),
      1927 => to_slv(opcode_type, 16#08#),
      1928 => to_slv(opcode_type, 16#09#),
      1929 => to_slv(opcode_type, 16#0E#),
      1930 => to_slv(opcode_type, 16#10#),
      1931 => to_slv(opcode_type, 16#07#),
      1932 => to_slv(opcode_type, 16#8D#),
      1933 => to_slv(opcode_type, 16#11#),
      1934 => to_slv(opcode_type, 16#07#),
      1935 => to_slv(opcode_type, 16#09#),
      1936 => to_slv(opcode_type, 16#0A#),
      1937 => to_slv(opcode_type, 16#10#),
      1938 => to_slv(opcode_type, 16#06#),
      1939 => to_slv(opcode_type, 16#10#),
      1940 => to_slv(opcode_type, 16#0E#),
      1941 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#07#),
      1953 => to_slv(opcode_type, 16#04#),
      1954 => to_slv(opcode_type, 16#01#),
      1955 => to_slv(opcode_type, 16#08#),
      1956 => to_slv(opcode_type, 16#0A#),
      1957 => to_slv(opcode_type, 16#0D#),
      1958 => to_slv(opcode_type, 16#09#),
      1959 => to_slv(opcode_type, 16#07#),
      1960 => to_slv(opcode_type, 16#06#),
      1961 => to_slv(opcode_type, 16#0F#),
      1962 => to_slv(opcode_type, 16#0D#),
      1963 => to_slv(opcode_type, 16#07#),
      1964 => to_slv(opcode_type, 16#BB#),
      1965 => to_slv(opcode_type, 16#0D#),
      1966 => to_slv(opcode_type, 16#09#),
      1967 => to_slv(opcode_type, 16#06#),
      1968 => to_slv(opcode_type, 16#16#),
      1969 => to_slv(opcode_type, 16#0C#),
      1970 => to_slv(opcode_type, 16#07#),
      1971 => to_slv(opcode_type, 16#11#),
      1972 => to_slv(opcode_type, 16#0B#),
      1973 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#07#),
      1985 => to_slv(opcode_type, 16#07#),
      1986 => to_slv(opcode_type, 16#01#),
      1987 => to_slv(opcode_type, 16#08#),
      1988 => to_slv(opcode_type, 16#0C#),
      1989 => to_slv(opcode_type, 16#93#),
      1990 => to_slv(opcode_type, 16#05#),
      1991 => to_slv(opcode_type, 16#07#),
      1992 => to_slv(opcode_type, 16#90#),
      1993 => to_slv(opcode_type, 16#0F#),
      1994 => to_slv(opcode_type, 16#07#),
      1995 => to_slv(opcode_type, 16#01#),
      1996 => to_slv(opcode_type, 16#04#),
      1997 => to_slv(opcode_type, 16#0B#),
      1998 => to_slv(opcode_type, 16#08#),
      1999 => to_slv(opcode_type, 16#09#),
      2000 => to_slv(opcode_type, 16#0E#),
      2001 => to_slv(opcode_type, 16#B7#),
      2002 => to_slv(opcode_type, 16#08#),
      2003 => to_slv(opcode_type, 16#0A#),
      2004 => to_slv(opcode_type, 16#0A#),
      2005 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#07#),
      2017 => to_slv(opcode_type, 16#04#),
      2018 => to_slv(opcode_type, 16#08#),
      2019 => to_slv(opcode_type, 16#06#),
      2020 => to_slv(opcode_type, 16#D8#),
      2021 => to_slv(opcode_type, 16#10#),
      2022 => to_slv(opcode_type, 16#07#),
      2023 => to_slv(opcode_type, 16#10#),
      2024 => to_slv(opcode_type, 16#0B#),
      2025 => to_slv(opcode_type, 16#06#),
      2026 => to_slv(opcode_type, 16#09#),
      2027 => to_slv(opcode_type, 16#06#),
      2028 => to_slv(opcode_type, 16#0F#),
      2029 => to_slv(opcode_type, 16#0A#),
      2030 => to_slv(opcode_type, 16#05#),
      2031 => to_slv(opcode_type, 16#0B#),
      2032 => to_slv(opcode_type, 16#06#),
      2033 => to_slv(opcode_type, 16#03#),
      2034 => to_slv(opcode_type, 16#10#),
      2035 => to_slv(opcode_type, 16#03#),
      2036 => to_slv(opcode_type, 16#0A#),
      2037 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#09#),
      2049 => to_slv(opcode_type, 16#06#),
      2050 => to_slv(opcode_type, 16#05#),
      2051 => to_slv(opcode_type, 16#08#),
      2052 => to_slv(opcode_type, 16#0D#),
      2053 => to_slv(opcode_type, 16#AB#),
      2054 => to_slv(opcode_type, 16#03#),
      2055 => to_slv(opcode_type, 16#03#),
      2056 => to_slv(opcode_type, 16#0B#),
      2057 => to_slv(opcode_type, 16#08#),
      2058 => to_slv(opcode_type, 16#03#),
      2059 => to_slv(opcode_type, 16#07#),
      2060 => to_slv(opcode_type, 16#0C#),
      2061 => to_slv(opcode_type, 16#0D#),
      2062 => to_slv(opcode_type, 16#08#),
      2063 => to_slv(opcode_type, 16#09#),
      2064 => to_slv(opcode_type, 16#0E#),
      2065 => to_slv(opcode_type, 16#0A#),
      2066 => to_slv(opcode_type, 16#08#),
      2067 => to_slv(opcode_type, 16#0A#),
      2068 => to_slv(opcode_type, 16#82#),
      2069 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#08#),
      2081 => to_slv(opcode_type, 16#01#),
      2082 => to_slv(opcode_type, 16#04#),
      2083 => to_slv(opcode_type, 16#08#),
      2084 => to_slv(opcode_type, 16#BD#),
      2085 => to_slv(opcode_type, 16#11#),
      2086 => to_slv(opcode_type, 16#09#),
      2087 => to_slv(opcode_type, 16#06#),
      2088 => to_slv(opcode_type, 16#07#),
      2089 => to_slv(opcode_type, 16#0C#),
      2090 => to_slv(opcode_type, 16#13#),
      2091 => to_slv(opcode_type, 16#08#),
      2092 => to_slv(opcode_type, 16#0F#),
      2093 => to_slv(opcode_type, 16#26#),
      2094 => to_slv(opcode_type, 16#08#),
      2095 => to_slv(opcode_type, 16#07#),
      2096 => to_slv(opcode_type, 16#63#),
      2097 => to_slv(opcode_type, 16#C7#),
      2098 => to_slv(opcode_type, 16#07#),
      2099 => to_slv(opcode_type, 16#0E#),
      2100 => to_slv(opcode_type, 16#0D#),
      2101 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#06#),
      2113 => to_slv(opcode_type, 16#01#),
      2114 => to_slv(opcode_type, 16#06#),
      2115 => to_slv(opcode_type, 16#05#),
      2116 => to_slv(opcode_type, 16#0D#),
      2117 => to_slv(opcode_type, 16#05#),
      2118 => to_slv(opcode_type, 16#0D#),
      2119 => to_slv(opcode_type, 16#07#),
      2120 => to_slv(opcode_type, 16#07#),
      2121 => to_slv(opcode_type, 16#08#),
      2122 => to_slv(opcode_type, 16#11#),
      2123 => to_slv(opcode_type, 16#0F#),
      2124 => to_slv(opcode_type, 16#05#),
      2125 => to_slv(opcode_type, 16#0D#),
      2126 => to_slv(opcode_type, 16#06#),
      2127 => to_slv(opcode_type, 16#06#),
      2128 => to_slv(opcode_type, 16#0F#),
      2129 => to_slv(opcode_type, 16#0E#),
      2130 => to_slv(opcode_type, 16#08#),
      2131 => to_slv(opcode_type, 16#33#),
      2132 => to_slv(opcode_type, 16#0A#),
      2133 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#09#),
      2146 => to_slv(opcode_type, 16#09#),
      2147 => to_slv(opcode_type, 16#04#),
      2148 => to_slv(opcode_type, 16#0C#),
      2149 => to_slv(opcode_type, 16#03#),
      2150 => to_slv(opcode_type, 16#0C#),
      2151 => to_slv(opcode_type, 16#05#),
      2152 => to_slv(opcode_type, 16#02#),
      2153 => to_slv(opcode_type, 16#11#),
      2154 => to_slv(opcode_type, 16#08#),
      2155 => to_slv(opcode_type, 16#08#),
      2156 => to_slv(opcode_type, 16#08#),
      2157 => to_slv(opcode_type, 16#0B#),
      2158 => to_slv(opcode_type, 16#0E#),
      2159 => to_slv(opcode_type, 16#07#),
      2160 => to_slv(opcode_type, 16#11#),
      2161 => to_slv(opcode_type, 16#0E#),
      2162 => to_slv(opcode_type, 16#04#),
      2163 => to_slv(opcode_type, 16#02#),
      2164 => to_slv(opcode_type, 16#0C#),
      2165 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#06#),
      2177 => to_slv(opcode_type, 16#05#),
      2178 => to_slv(opcode_type, 16#05#),
      2179 => to_slv(opcode_type, 16#07#),
      2180 => to_slv(opcode_type, 16#0D#),
      2181 => to_slv(opcode_type, 16#0F#),
      2182 => to_slv(opcode_type, 16#09#),
      2183 => to_slv(opcode_type, 16#06#),
      2184 => to_slv(opcode_type, 16#06#),
      2185 => to_slv(opcode_type, 16#F0#),
      2186 => to_slv(opcode_type, 16#0B#),
      2187 => to_slv(opcode_type, 16#08#),
      2188 => to_slv(opcode_type, 16#0C#),
      2189 => to_slv(opcode_type, 16#0C#),
      2190 => to_slv(opcode_type, 16#07#),
      2191 => to_slv(opcode_type, 16#09#),
      2192 => to_slv(opcode_type, 16#0E#),
      2193 => to_slv(opcode_type, 16#0B#),
      2194 => to_slv(opcode_type, 16#06#),
      2195 => to_slv(opcode_type, 16#30#),
      2196 => to_slv(opcode_type, 16#0A#),
      2197 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#08#),
      2209 => to_slv(opcode_type, 16#05#),
      2210 => to_slv(opcode_type, 16#06#),
      2211 => to_slv(opcode_type, 16#04#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#07#),
      2214 => to_slv(opcode_type, 16#0E#),
      2215 => to_slv(opcode_type, 16#10#),
      2216 => to_slv(opcode_type, 16#09#),
      2217 => to_slv(opcode_type, 16#06#),
      2218 => to_slv(opcode_type, 16#03#),
      2219 => to_slv(opcode_type, 16#0C#),
      2220 => to_slv(opcode_type, 16#08#),
      2221 => to_slv(opcode_type, 16#11#),
      2222 => to_slv(opcode_type, 16#0C#),
      2223 => to_slv(opcode_type, 16#07#),
      2224 => to_slv(opcode_type, 16#05#),
      2225 => to_slv(opcode_type, 16#0F#),
      2226 => to_slv(opcode_type, 16#07#),
      2227 => to_slv(opcode_type, 16#0C#),
      2228 => to_slv(opcode_type, 16#0C#),
      2229 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#09#),
      2241 => to_slv(opcode_type, 16#06#),
      2242 => to_slv(opcode_type, 16#01#),
      2243 => to_slv(opcode_type, 16#01#),
      2244 => to_slv(opcode_type, 16#0B#),
      2245 => to_slv(opcode_type, 16#02#),
      2246 => to_slv(opcode_type, 16#09#),
      2247 => to_slv(opcode_type, 16#0F#),
      2248 => to_slv(opcode_type, 16#11#),
      2249 => to_slv(opcode_type, 16#07#),
      2250 => to_slv(opcode_type, 16#03#),
      2251 => to_slv(opcode_type, 16#07#),
      2252 => to_slv(opcode_type, 16#0A#),
      2253 => to_slv(opcode_type, 16#0D#),
      2254 => to_slv(opcode_type, 16#07#),
      2255 => to_slv(opcode_type, 16#08#),
      2256 => to_slv(opcode_type, 16#0E#),
      2257 => to_slv(opcode_type, 16#0E#),
      2258 => to_slv(opcode_type, 16#07#),
      2259 => to_slv(opcode_type, 16#0F#),
      2260 => to_slv(opcode_type, 16#0A#),
      2261 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#07#),
      2273 => to_slv(opcode_type, 16#03#),
      2274 => to_slv(opcode_type, 16#07#),
      2275 => to_slv(opcode_type, 16#02#),
      2276 => to_slv(opcode_type, 16#10#),
      2277 => to_slv(opcode_type, 16#07#),
      2278 => to_slv(opcode_type, 16#10#),
      2279 => to_slv(opcode_type, 16#0A#),
      2280 => to_slv(opcode_type, 16#08#),
      2281 => to_slv(opcode_type, 16#08#),
      2282 => to_slv(opcode_type, 16#09#),
      2283 => to_slv(opcode_type, 16#0C#),
      2284 => to_slv(opcode_type, 16#0D#),
      2285 => to_slv(opcode_type, 16#02#),
      2286 => to_slv(opcode_type, 16#10#),
      2287 => to_slv(opcode_type, 16#09#),
      2288 => to_slv(opcode_type, 16#03#),
      2289 => to_slv(opcode_type, 16#11#),
      2290 => to_slv(opcode_type, 16#07#),
      2291 => to_slv(opcode_type, 16#0A#),
      2292 => to_slv(opcode_type, 16#11#),
      2293 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#08#),
      2305 => to_slv(opcode_type, 16#05#),
      2306 => to_slv(opcode_type, 16#07#),
      2307 => to_slv(opcode_type, 16#04#),
      2308 => to_slv(opcode_type, 16#0D#),
      2309 => to_slv(opcode_type, 16#09#),
      2310 => to_slv(opcode_type, 16#0F#),
      2311 => to_slv(opcode_type, 16#0B#),
      2312 => to_slv(opcode_type, 16#09#),
      2313 => to_slv(opcode_type, 16#06#),
      2314 => to_slv(opcode_type, 16#08#),
      2315 => to_slv(opcode_type, 16#0C#),
      2316 => to_slv(opcode_type, 16#10#),
      2317 => to_slv(opcode_type, 16#04#),
      2318 => to_slv(opcode_type, 16#0B#),
      2319 => to_slv(opcode_type, 16#06#),
      2320 => to_slv(opcode_type, 16#02#),
      2321 => to_slv(opcode_type, 16#0B#),
      2322 => to_slv(opcode_type, 16#06#),
      2323 => to_slv(opcode_type, 16#0A#),
      2324 => to_slv(opcode_type, 16#0A#),
      2325 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#08#),
      2337 => to_slv(opcode_type, 16#07#),
      2338 => to_slv(opcode_type, 16#03#),
      2339 => to_slv(opcode_type, 16#01#),
      2340 => to_slv(opcode_type, 16#0B#),
      2341 => to_slv(opcode_type, 16#09#),
      2342 => to_slv(opcode_type, 16#05#),
      2343 => to_slv(opcode_type, 16#30#),
      2344 => to_slv(opcode_type, 16#09#),
      2345 => to_slv(opcode_type, 16#0E#),
      2346 => to_slv(opcode_type, 16#0F#),
      2347 => to_slv(opcode_type, 16#09#),
      2348 => to_slv(opcode_type, 16#03#),
      2349 => to_slv(opcode_type, 16#08#),
      2350 => to_slv(opcode_type, 16#0E#),
      2351 => to_slv(opcode_type, 16#0D#),
      2352 => to_slv(opcode_type, 16#08#),
      2353 => to_slv(opcode_type, 16#06#),
      2354 => to_slv(opcode_type, 16#0F#),
      2355 => to_slv(opcode_type, 16#0C#),
      2356 => to_slv(opcode_type, 16#0C#),
      2357 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#08#),
      2369 => to_slv(opcode_type, 16#05#),
      2370 => to_slv(opcode_type, 16#02#),
      2371 => to_slv(opcode_type, 16#07#),
      2372 => to_slv(opcode_type, 16#0D#),
      2373 => to_slv(opcode_type, 16#0B#),
      2374 => to_slv(opcode_type, 16#07#),
      2375 => to_slv(opcode_type, 16#06#),
      2376 => to_slv(opcode_type, 16#07#),
      2377 => to_slv(opcode_type, 16#0C#),
      2378 => to_slv(opcode_type, 16#0B#),
      2379 => to_slv(opcode_type, 16#07#),
      2380 => to_slv(opcode_type, 16#0C#),
      2381 => to_slv(opcode_type, 16#0C#),
      2382 => to_slv(opcode_type, 16#09#),
      2383 => to_slv(opcode_type, 16#08#),
      2384 => to_slv(opcode_type, 16#0D#),
      2385 => to_slv(opcode_type, 16#0B#),
      2386 => to_slv(opcode_type, 16#06#),
      2387 => to_slv(opcode_type, 16#0D#),
      2388 => to_slv(opcode_type, 16#10#),
      2389 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#08#),
      2402 => to_slv(opcode_type, 16#04#),
      2403 => to_slv(opcode_type, 16#05#),
      2404 => to_slv(opcode_type, 16#10#),
      2405 => to_slv(opcode_type, 16#09#),
      2406 => to_slv(opcode_type, 16#03#),
      2407 => to_slv(opcode_type, 16#0E#),
      2408 => to_slv(opcode_type, 16#08#),
      2409 => to_slv(opcode_type, 16#0D#),
      2410 => to_slv(opcode_type, 16#0F#),
      2411 => to_slv(opcode_type, 16#07#),
      2412 => to_slv(opcode_type, 16#01#),
      2413 => to_slv(opcode_type, 16#01#),
      2414 => to_slv(opcode_type, 16#59#),
      2415 => to_slv(opcode_type, 16#06#),
      2416 => to_slv(opcode_type, 16#04#),
      2417 => to_slv(opcode_type, 16#11#),
      2418 => to_slv(opcode_type, 16#08#),
      2419 => to_slv(opcode_type, 16#0B#),
      2420 => to_slv(opcode_type, 16#0D#),
      2421 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#09#),
      2433 => to_slv(opcode_type, 16#05#),
      2434 => to_slv(opcode_type, 16#06#),
      2435 => to_slv(opcode_type, 16#07#),
      2436 => to_slv(opcode_type, 16#0A#),
      2437 => to_slv(opcode_type, 16#10#),
      2438 => to_slv(opcode_type, 16#06#),
      2439 => to_slv(opcode_type, 16#3F#),
      2440 => to_slv(opcode_type, 16#41#),
      2441 => to_slv(opcode_type, 16#06#),
      2442 => to_slv(opcode_type, 16#03#),
      2443 => to_slv(opcode_type, 16#06#),
      2444 => to_slv(opcode_type, 16#0E#),
      2445 => to_slv(opcode_type, 16#0B#),
      2446 => to_slv(opcode_type, 16#06#),
      2447 => to_slv(opcode_type, 16#08#),
      2448 => to_slv(opcode_type, 16#1A#),
      2449 => to_slv(opcode_type, 16#11#),
      2450 => to_slv(opcode_type, 16#06#),
      2451 => to_slv(opcode_type, 16#0B#),
      2452 => to_slv(opcode_type, 16#0C#),
      2453 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#08#),
      2465 => to_slv(opcode_type, 16#09#),
      2466 => to_slv(opcode_type, 16#07#),
      2467 => to_slv(opcode_type, 16#05#),
      2468 => to_slv(opcode_type, 16#52#),
      2469 => to_slv(opcode_type, 16#02#),
      2470 => to_slv(opcode_type, 16#0C#),
      2471 => to_slv(opcode_type, 16#06#),
      2472 => to_slv(opcode_type, 16#09#),
      2473 => to_slv(opcode_type, 16#0A#),
      2474 => to_slv(opcode_type, 16#0D#),
      2475 => to_slv(opcode_type, 16#09#),
      2476 => to_slv(opcode_type, 16#0C#),
      2477 => to_slv(opcode_type, 16#0D#),
      2478 => to_slv(opcode_type, 16#04#),
      2479 => to_slv(opcode_type, 16#07#),
      2480 => to_slv(opcode_type, 16#06#),
      2481 => to_slv(opcode_type, 16#0F#),
      2482 => to_slv(opcode_type, 16#0E#),
      2483 => to_slv(opcode_type, 16#05#),
      2484 => to_slv(opcode_type, 16#0A#),
      2485 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#07#),
      2497 => to_slv(opcode_type, 16#09#),
      2498 => to_slv(opcode_type, 16#06#),
      2499 => to_slv(opcode_type, 16#09#),
      2500 => to_slv(opcode_type, 16#0B#),
      2501 => to_slv(opcode_type, 16#0F#),
      2502 => to_slv(opcode_type, 16#08#),
      2503 => to_slv(opcode_type, 16#0F#),
      2504 => to_slv(opcode_type, 16#10#),
      2505 => to_slv(opcode_type, 16#07#),
      2506 => to_slv(opcode_type, 16#08#),
      2507 => to_slv(opcode_type, 16#0B#),
      2508 => to_slv(opcode_type, 16#0B#),
      2509 => to_slv(opcode_type, 16#03#),
      2510 => to_slv(opcode_type, 16#0E#),
      2511 => to_slv(opcode_type, 16#06#),
      2512 => to_slv(opcode_type, 16#03#),
      2513 => to_slv(opcode_type, 16#08#),
      2514 => to_slv(opcode_type, 16#0A#),
      2515 => to_slv(opcode_type, 16#0E#),
      2516 => to_slv(opcode_type, 16#0B#),
      2517 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#02#),
      2530 => to_slv(opcode_type, 16#01#),
      2531 => to_slv(opcode_type, 16#07#),
      2532 => to_slv(opcode_type, 16#0A#),
      2533 => to_slv(opcode_type, 16#0B#),
      2534 => to_slv(opcode_type, 16#08#),
      2535 => to_slv(opcode_type, 16#06#),
      2536 => to_slv(opcode_type, 16#06#),
      2537 => to_slv(opcode_type, 16#11#),
      2538 => to_slv(opcode_type, 16#0F#),
      2539 => to_slv(opcode_type, 16#09#),
      2540 => to_slv(opcode_type, 16#11#),
      2541 => to_slv(opcode_type, 16#0B#),
      2542 => to_slv(opcode_type, 16#06#),
      2543 => to_slv(opcode_type, 16#09#),
      2544 => to_slv(opcode_type, 16#C2#),
      2545 => to_slv(opcode_type, 16#10#),
      2546 => to_slv(opcode_type, 16#07#),
      2547 => to_slv(opcode_type, 16#0C#),
      2548 => to_slv(opcode_type, 16#0E#),
      2549 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#09#),
      2561 => to_slv(opcode_type, 16#03#),
      2562 => to_slv(opcode_type, 16#02#),
      2563 => to_slv(opcode_type, 16#08#),
      2564 => to_slv(opcode_type, 16#0E#),
      2565 => to_slv(opcode_type, 16#0D#),
      2566 => to_slv(opcode_type, 16#06#),
      2567 => to_slv(opcode_type, 16#07#),
      2568 => to_slv(opcode_type, 16#07#),
      2569 => to_slv(opcode_type, 16#10#),
      2570 => to_slv(opcode_type, 16#7F#),
      2571 => to_slv(opcode_type, 16#09#),
      2572 => to_slv(opcode_type, 16#0A#),
      2573 => to_slv(opcode_type, 16#11#),
      2574 => to_slv(opcode_type, 16#09#),
      2575 => to_slv(opcode_type, 16#07#),
      2576 => to_slv(opcode_type, 16#11#),
      2577 => to_slv(opcode_type, 16#0D#),
      2578 => to_slv(opcode_type, 16#09#),
      2579 => to_slv(opcode_type, 16#10#),
      2580 => to_slv(opcode_type, 16#0E#),
      2581 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#06#),
      2593 => to_slv(opcode_type, 16#09#),
      2594 => to_slv(opcode_type, 16#06#),
      2595 => to_slv(opcode_type, 16#07#),
      2596 => to_slv(opcode_type, 16#0C#),
      2597 => to_slv(opcode_type, 16#0F#),
      2598 => to_slv(opcode_type, 16#05#),
      2599 => to_slv(opcode_type, 16#0C#),
      2600 => to_slv(opcode_type, 16#09#),
      2601 => to_slv(opcode_type, 16#04#),
      2602 => to_slv(opcode_type, 16#10#),
      2603 => to_slv(opcode_type, 16#04#),
      2604 => to_slv(opcode_type, 16#11#),
      2605 => to_slv(opcode_type, 16#07#),
      2606 => to_slv(opcode_type, 16#05#),
      2607 => to_slv(opcode_type, 16#06#),
      2608 => to_slv(opcode_type, 16#0C#),
      2609 => to_slv(opcode_type, 16#0C#),
      2610 => to_slv(opcode_type, 16#08#),
      2611 => to_slv(opcode_type, 16#0B#),
      2612 => to_slv(opcode_type, 16#0D#),
      2613 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#08#),
      2625 => to_slv(opcode_type, 16#02#),
      2626 => to_slv(opcode_type, 16#05#),
      2627 => to_slv(opcode_type, 16#09#),
      2628 => to_slv(opcode_type, 16#0E#),
      2629 => to_slv(opcode_type, 16#11#),
      2630 => to_slv(opcode_type, 16#09#),
      2631 => to_slv(opcode_type, 16#08#),
      2632 => to_slv(opcode_type, 16#06#),
      2633 => to_slv(opcode_type, 16#0B#),
      2634 => to_slv(opcode_type, 16#0F#),
      2635 => to_slv(opcode_type, 16#07#),
      2636 => to_slv(opcode_type, 16#0F#),
      2637 => to_slv(opcode_type, 16#11#),
      2638 => to_slv(opcode_type, 16#07#),
      2639 => to_slv(opcode_type, 16#06#),
      2640 => to_slv(opcode_type, 16#0A#),
      2641 => to_slv(opcode_type, 16#10#),
      2642 => to_slv(opcode_type, 16#08#),
      2643 => to_slv(opcode_type, 16#0F#),
      2644 => to_slv(opcode_type, 16#CA#),
      2645 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#09#),
      2657 => to_slv(opcode_type, 16#09#),
      2658 => to_slv(opcode_type, 16#06#),
      2659 => to_slv(opcode_type, 16#04#),
      2660 => to_slv(opcode_type, 16#0A#),
      2661 => to_slv(opcode_type, 16#08#),
      2662 => to_slv(opcode_type, 16#10#),
      2663 => to_slv(opcode_type, 16#0F#),
      2664 => to_slv(opcode_type, 16#03#),
      2665 => to_slv(opcode_type, 16#07#),
      2666 => to_slv(opcode_type, 16#0F#),
      2667 => to_slv(opcode_type, 16#10#),
      2668 => to_slv(opcode_type, 16#09#),
      2669 => to_slv(opcode_type, 16#01#),
      2670 => to_slv(opcode_type, 16#01#),
      2671 => to_slv(opcode_type, 16#0D#),
      2672 => to_slv(opcode_type, 16#06#),
      2673 => to_slv(opcode_type, 16#09#),
      2674 => to_slv(opcode_type, 16#F6#),
      2675 => to_slv(opcode_type, 16#0D#),
      2676 => to_slv(opcode_type, 16#10#),
      2677 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#07#),
      2689 => to_slv(opcode_type, 16#06#),
      2690 => to_slv(opcode_type, 16#05#),
      2691 => to_slv(opcode_type, 16#02#),
      2692 => to_slv(opcode_type, 16#75#),
      2693 => to_slv(opcode_type, 16#08#),
      2694 => to_slv(opcode_type, 16#05#),
      2695 => to_slv(opcode_type, 16#0F#),
      2696 => to_slv(opcode_type, 16#06#),
      2697 => to_slv(opcode_type, 16#0D#),
      2698 => to_slv(opcode_type, 16#0B#),
      2699 => to_slv(opcode_type, 16#06#),
      2700 => to_slv(opcode_type, 16#09#),
      2701 => to_slv(opcode_type, 16#03#),
      2702 => to_slv(opcode_type, 16#19#),
      2703 => to_slv(opcode_type, 16#08#),
      2704 => to_slv(opcode_type, 16#66#),
      2705 => to_slv(opcode_type, 16#9D#),
      2706 => to_slv(opcode_type, 16#05#),
      2707 => to_slv(opcode_type, 16#04#),
      2708 => to_slv(opcode_type, 16#EF#),
      2709 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#09#),
      2721 => to_slv(opcode_type, 16#08#),
      2722 => to_slv(opcode_type, 16#07#),
      2723 => to_slv(opcode_type, 16#08#),
      2724 => to_slv(opcode_type, 16#0A#),
      2725 => to_slv(opcode_type, 16#0D#),
      2726 => to_slv(opcode_type, 16#02#),
      2727 => to_slv(opcode_type, 16#0D#),
      2728 => to_slv(opcode_type, 16#08#),
      2729 => to_slv(opcode_type, 16#09#),
      2730 => to_slv(opcode_type, 16#0C#),
      2731 => to_slv(opcode_type, 16#0B#),
      2732 => to_slv(opcode_type, 16#03#),
      2733 => to_slv(opcode_type, 16#CD#),
      2734 => to_slv(opcode_type, 16#02#),
      2735 => to_slv(opcode_type, 16#06#),
      2736 => to_slv(opcode_type, 16#04#),
      2737 => to_slv(opcode_type, 16#0C#),
      2738 => to_slv(opcode_type, 16#07#),
      2739 => to_slv(opcode_type, 16#11#),
      2740 => to_slv(opcode_type, 16#10#),
      2741 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#06#),
      2753 => to_slv(opcode_type, 16#05#),
      2754 => to_slv(opcode_type, 16#05#),
      2755 => to_slv(opcode_type, 16#08#),
      2756 => to_slv(opcode_type, 16#0D#),
      2757 => to_slv(opcode_type, 16#0D#),
      2758 => to_slv(opcode_type, 16#09#),
      2759 => to_slv(opcode_type, 16#09#),
      2760 => to_slv(opcode_type, 16#07#),
      2761 => to_slv(opcode_type, 16#0F#),
      2762 => to_slv(opcode_type, 16#10#),
      2763 => to_slv(opcode_type, 16#09#),
      2764 => to_slv(opcode_type, 16#0B#),
      2765 => to_slv(opcode_type, 16#0F#),
      2766 => to_slv(opcode_type, 16#07#),
      2767 => to_slv(opcode_type, 16#06#),
      2768 => to_slv(opcode_type, 16#0F#),
      2769 => to_slv(opcode_type, 16#B6#),
      2770 => to_slv(opcode_type, 16#07#),
      2771 => to_slv(opcode_type, 16#0E#),
      2772 => to_slv(opcode_type, 16#0B#),
      2773 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#06#),
      2785 => to_slv(opcode_type, 16#06#),
      2786 => to_slv(opcode_type, 16#09#),
      2787 => to_slv(opcode_type, 16#08#),
      2788 => to_slv(opcode_type, 16#10#),
      2789 => to_slv(opcode_type, 16#0D#),
      2790 => to_slv(opcode_type, 16#05#),
      2791 => to_slv(opcode_type, 16#0F#),
      2792 => to_slv(opcode_type, 16#06#),
      2793 => to_slv(opcode_type, 16#01#),
      2794 => to_slv(opcode_type, 16#0A#),
      2795 => to_slv(opcode_type, 16#01#),
      2796 => to_slv(opcode_type, 16#0B#),
      2797 => to_slv(opcode_type, 16#03#),
      2798 => to_slv(opcode_type, 16#09#),
      2799 => to_slv(opcode_type, 16#08#),
      2800 => to_slv(opcode_type, 16#B7#),
      2801 => to_slv(opcode_type, 16#0A#),
      2802 => to_slv(opcode_type, 16#07#),
      2803 => to_slv(opcode_type, 16#0B#),
      2804 => to_slv(opcode_type, 16#10#),
      2805 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#07#),
      2817 => to_slv(opcode_type, 16#05#),
      2818 => to_slv(opcode_type, 16#02#),
      2819 => to_slv(opcode_type, 16#08#),
      2820 => to_slv(opcode_type, 16#0F#),
      2821 => to_slv(opcode_type, 16#0F#),
      2822 => to_slv(opcode_type, 16#06#),
      2823 => to_slv(opcode_type, 16#09#),
      2824 => to_slv(opcode_type, 16#08#),
      2825 => to_slv(opcode_type, 16#0A#),
      2826 => to_slv(opcode_type, 16#0C#),
      2827 => to_slv(opcode_type, 16#09#),
      2828 => to_slv(opcode_type, 16#0E#),
      2829 => to_slv(opcode_type, 16#0F#),
      2830 => to_slv(opcode_type, 16#09#),
      2831 => to_slv(opcode_type, 16#09#),
      2832 => to_slv(opcode_type, 16#0D#),
      2833 => to_slv(opcode_type, 16#0D#),
      2834 => to_slv(opcode_type, 16#07#),
      2835 => to_slv(opcode_type, 16#6C#),
      2836 => to_slv(opcode_type, 16#0F#),
      2837 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#09#),
      2849 => to_slv(opcode_type, 16#07#),
      2850 => to_slv(opcode_type, 16#07#),
      2851 => to_slv(opcode_type, 16#06#),
      2852 => to_slv(opcode_type, 16#11#),
      2853 => to_slv(opcode_type, 16#0F#),
      2854 => to_slv(opcode_type, 16#09#),
      2855 => to_slv(opcode_type, 16#BA#),
      2856 => to_slv(opcode_type, 16#0D#),
      2857 => to_slv(opcode_type, 16#08#),
      2858 => to_slv(opcode_type, 16#05#),
      2859 => to_slv(opcode_type, 16#0A#),
      2860 => to_slv(opcode_type, 16#04#),
      2861 => to_slv(opcode_type, 16#0F#),
      2862 => to_slv(opcode_type, 16#06#),
      2863 => to_slv(opcode_type, 16#05#),
      2864 => to_slv(opcode_type, 16#03#),
      2865 => to_slv(opcode_type, 16#0F#),
      2866 => to_slv(opcode_type, 16#06#),
      2867 => to_slv(opcode_type, 16#0C#),
      2868 => to_slv(opcode_type, 16#0D#),
      2869 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#07#),
      2881 => to_slv(opcode_type, 16#02#),
      2882 => to_slv(opcode_type, 16#02#),
      2883 => to_slv(opcode_type, 16#08#),
      2884 => to_slv(opcode_type, 16#0C#),
      2885 => to_slv(opcode_type, 16#5D#),
      2886 => to_slv(opcode_type, 16#09#),
      2887 => to_slv(opcode_type, 16#09#),
      2888 => to_slv(opcode_type, 16#06#),
      2889 => to_slv(opcode_type, 16#0A#),
      2890 => to_slv(opcode_type, 16#11#),
      2891 => to_slv(opcode_type, 16#07#),
      2892 => to_slv(opcode_type, 16#11#),
      2893 => to_slv(opcode_type, 16#27#),
      2894 => to_slv(opcode_type, 16#06#),
      2895 => to_slv(opcode_type, 16#06#),
      2896 => to_slv(opcode_type, 16#2B#),
      2897 => to_slv(opcode_type, 16#78#),
      2898 => to_slv(opcode_type, 16#09#),
      2899 => to_slv(opcode_type, 16#0D#),
      2900 => to_slv(opcode_type, 16#A2#),
      2901 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#07#),
      2913 => to_slv(opcode_type, 16#05#),
      2914 => to_slv(opcode_type, 16#07#),
      2915 => to_slv(opcode_type, 16#08#),
      2916 => to_slv(opcode_type, 16#8A#),
      2917 => to_slv(opcode_type, 16#0F#),
      2918 => to_slv(opcode_type, 16#06#),
      2919 => to_slv(opcode_type, 16#0F#),
      2920 => to_slv(opcode_type, 16#0A#),
      2921 => to_slv(opcode_type, 16#09#),
      2922 => to_slv(opcode_type, 16#07#),
      2923 => to_slv(opcode_type, 16#09#),
      2924 => to_slv(opcode_type, 16#0C#),
      2925 => to_slv(opcode_type, 16#0F#),
      2926 => to_slv(opcode_type, 16#02#),
      2927 => to_slv(opcode_type, 16#0C#),
      2928 => to_slv(opcode_type, 16#07#),
      2929 => to_slv(opcode_type, 16#02#),
      2930 => to_slv(opcode_type, 16#11#),
      2931 => to_slv(opcode_type, 16#05#),
      2932 => to_slv(opcode_type, 16#0B#),
      2933 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#08#),
      2945 => to_slv(opcode_type, 16#05#),
      2946 => to_slv(opcode_type, 16#02#),
      2947 => to_slv(opcode_type, 16#09#),
      2948 => to_slv(opcode_type, 16#0B#),
      2949 => to_slv(opcode_type, 16#11#),
      2950 => to_slv(opcode_type, 16#09#),
      2951 => to_slv(opcode_type, 16#09#),
      2952 => to_slv(opcode_type, 16#06#),
      2953 => to_slv(opcode_type, 16#0E#),
      2954 => to_slv(opcode_type, 16#10#),
      2955 => to_slv(opcode_type, 16#06#),
      2956 => to_slv(opcode_type, 16#28#),
      2957 => to_slv(opcode_type, 16#0F#),
      2958 => to_slv(opcode_type, 16#09#),
      2959 => to_slv(opcode_type, 16#07#),
      2960 => to_slv(opcode_type, 16#0B#),
      2961 => to_slv(opcode_type, 16#0A#),
      2962 => to_slv(opcode_type, 16#06#),
      2963 => to_slv(opcode_type, 16#0C#),
      2964 => to_slv(opcode_type, 16#0D#),
      2965 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#09#),
      2977 => to_slv(opcode_type, 16#07#),
      2978 => to_slv(opcode_type, 16#06#),
      2979 => to_slv(opcode_type, 16#02#),
      2980 => to_slv(opcode_type, 16#0C#),
      2981 => to_slv(opcode_type, 16#06#),
      2982 => to_slv(opcode_type, 16#0A#),
      2983 => to_slv(opcode_type, 16#0D#),
      2984 => to_slv(opcode_type, 16#03#),
      2985 => to_slv(opcode_type, 16#03#),
      2986 => to_slv(opcode_type, 16#0D#),
      2987 => to_slv(opcode_type, 16#09#),
      2988 => to_slv(opcode_type, 16#02#),
      2989 => to_slv(opcode_type, 16#03#),
      2990 => to_slv(opcode_type, 16#0A#),
      2991 => to_slv(opcode_type, 16#08#),
      2992 => to_slv(opcode_type, 16#09#),
      2993 => to_slv(opcode_type, 16#11#),
      2994 => to_slv(opcode_type, 16#0F#),
      2995 => to_slv(opcode_type, 16#05#),
      2996 => to_slv(opcode_type, 16#0F#),
      2997 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#06#),
      3009 => to_slv(opcode_type, 16#03#),
      3010 => to_slv(opcode_type, 16#01#),
      3011 => to_slv(opcode_type, 16#06#),
      3012 => to_slv(opcode_type, 16#11#),
      3013 => to_slv(opcode_type, 16#0D#),
      3014 => to_slv(opcode_type, 16#08#),
      3015 => to_slv(opcode_type, 16#07#),
      3016 => to_slv(opcode_type, 16#08#),
      3017 => to_slv(opcode_type, 16#10#),
      3018 => to_slv(opcode_type, 16#0E#),
      3019 => to_slv(opcode_type, 16#09#),
      3020 => to_slv(opcode_type, 16#0D#),
      3021 => to_slv(opcode_type, 16#0A#),
      3022 => to_slv(opcode_type, 16#07#),
      3023 => to_slv(opcode_type, 16#09#),
      3024 => to_slv(opcode_type, 16#0E#),
      3025 => to_slv(opcode_type, 16#0A#),
      3026 => to_slv(opcode_type, 16#07#),
      3027 => to_slv(opcode_type, 16#11#),
      3028 => to_slv(opcode_type, 16#0D#),
      3029 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#07#),
      3041 => to_slv(opcode_type, 16#07#),
      3042 => to_slv(opcode_type, 16#08#),
      3043 => to_slv(opcode_type, 16#02#),
      3044 => to_slv(opcode_type, 16#0E#),
      3045 => to_slv(opcode_type, 16#09#),
      3046 => to_slv(opcode_type, 16#0B#),
      3047 => to_slv(opcode_type, 16#89#),
      3048 => to_slv(opcode_type, 16#07#),
      3049 => to_slv(opcode_type, 16#08#),
      3050 => to_slv(opcode_type, 16#0D#),
      3051 => to_slv(opcode_type, 16#10#),
      3052 => to_slv(opcode_type, 16#05#),
      3053 => to_slv(opcode_type, 16#0A#),
      3054 => to_slv(opcode_type, 16#06#),
      3055 => to_slv(opcode_type, 16#09#),
      3056 => to_slv(opcode_type, 16#03#),
      3057 => to_slv(opcode_type, 16#11#),
      3058 => to_slv(opcode_type, 16#02#),
      3059 => to_slv(opcode_type, 16#0D#),
      3060 => to_slv(opcode_type, 16#0F#),
      3061 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#08#),
      3073 => to_slv(opcode_type, 16#07#),
      3074 => to_slv(opcode_type, 16#04#),
      3075 => to_slv(opcode_type, 16#01#),
      3076 => to_slv(opcode_type, 16#0E#),
      3077 => to_slv(opcode_type, 16#02#),
      3078 => to_slv(opcode_type, 16#06#),
      3079 => to_slv(opcode_type, 16#0D#),
      3080 => to_slv(opcode_type, 16#0A#),
      3081 => to_slv(opcode_type, 16#09#),
      3082 => to_slv(opcode_type, 16#01#),
      3083 => to_slv(opcode_type, 16#06#),
      3084 => to_slv(opcode_type, 16#11#),
      3085 => to_slv(opcode_type, 16#0D#),
      3086 => to_slv(opcode_type, 16#06#),
      3087 => to_slv(opcode_type, 16#08#),
      3088 => to_slv(opcode_type, 16#11#),
      3089 => to_slv(opcode_type, 16#0D#),
      3090 => to_slv(opcode_type, 16#09#),
      3091 => to_slv(opcode_type, 16#0D#),
      3092 => to_slv(opcode_type, 16#D8#),
      3093 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#08#),
      3105 => to_slv(opcode_type, 16#02#),
      3106 => to_slv(opcode_type, 16#09#),
      3107 => to_slv(opcode_type, 16#01#),
      3108 => to_slv(opcode_type, 16#0B#),
      3109 => to_slv(opcode_type, 16#03#),
      3110 => to_slv(opcode_type, 16#0C#),
      3111 => to_slv(opcode_type, 16#07#),
      3112 => to_slv(opcode_type, 16#07#),
      3113 => to_slv(opcode_type, 16#06#),
      3114 => to_slv(opcode_type, 16#11#),
      3115 => to_slv(opcode_type, 16#0F#),
      3116 => to_slv(opcode_type, 16#03#),
      3117 => to_slv(opcode_type, 16#10#),
      3118 => to_slv(opcode_type, 16#06#),
      3119 => to_slv(opcode_type, 16#06#),
      3120 => to_slv(opcode_type, 16#0B#),
      3121 => to_slv(opcode_type, 16#0F#),
      3122 => to_slv(opcode_type, 16#08#),
      3123 => to_slv(opcode_type, 16#10#),
      3124 => to_slv(opcode_type, 16#11#),
      3125 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#09#),
      3137 => to_slv(opcode_type, 16#09#),
      3138 => to_slv(opcode_type, 16#04#),
      3139 => to_slv(opcode_type, 16#09#),
      3140 => to_slv(opcode_type, 16#10#),
      3141 => to_slv(opcode_type, 16#FC#),
      3142 => to_slv(opcode_type, 16#03#),
      3143 => to_slv(opcode_type, 16#09#),
      3144 => to_slv(opcode_type, 16#0E#),
      3145 => to_slv(opcode_type, 16#0B#),
      3146 => to_slv(opcode_type, 16#09#),
      3147 => to_slv(opcode_type, 16#04#),
      3148 => to_slv(opcode_type, 16#04#),
      3149 => to_slv(opcode_type, 16#0B#),
      3150 => to_slv(opcode_type, 16#08#),
      3151 => to_slv(opcode_type, 16#09#),
      3152 => to_slv(opcode_type, 16#0F#),
      3153 => to_slv(opcode_type, 16#0D#),
      3154 => to_slv(opcode_type, 16#06#),
      3155 => to_slv(opcode_type, 16#0E#),
      3156 => to_slv(opcode_type, 16#0C#),
      3157 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#06#),
      3169 => to_slv(opcode_type, 16#03#),
      3170 => to_slv(opcode_type, 16#05#),
      3171 => to_slv(opcode_type, 16#09#),
      3172 => to_slv(opcode_type, 16#0B#),
      3173 => to_slv(opcode_type, 16#0A#),
      3174 => to_slv(opcode_type, 16#09#),
      3175 => to_slv(opcode_type, 16#07#),
      3176 => to_slv(opcode_type, 16#09#),
      3177 => to_slv(opcode_type, 16#11#),
      3178 => to_slv(opcode_type, 16#0F#),
      3179 => to_slv(opcode_type, 16#06#),
      3180 => to_slv(opcode_type, 16#0C#),
      3181 => to_slv(opcode_type, 16#0A#),
      3182 => to_slv(opcode_type, 16#07#),
      3183 => to_slv(opcode_type, 16#06#),
      3184 => to_slv(opcode_type, 16#0E#),
      3185 => to_slv(opcode_type, 16#0F#),
      3186 => to_slv(opcode_type, 16#09#),
      3187 => to_slv(opcode_type, 16#0C#),
      3188 => to_slv(opcode_type, 16#0A#),
      3189 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#07#),
      3201 => to_slv(opcode_type, 16#07#),
      3202 => to_slv(opcode_type, 16#04#),
      3203 => to_slv(opcode_type, 16#03#),
      3204 => to_slv(opcode_type, 16#0F#),
      3205 => to_slv(opcode_type, 16#08#),
      3206 => to_slv(opcode_type, 16#09#),
      3207 => to_slv(opcode_type, 16#0C#),
      3208 => to_slv(opcode_type, 16#0F#),
      3209 => to_slv(opcode_type, 16#06#),
      3210 => to_slv(opcode_type, 16#10#),
      3211 => to_slv(opcode_type, 16#0B#),
      3212 => to_slv(opcode_type, 16#08#),
      3213 => to_slv(opcode_type, 16#04#),
      3214 => to_slv(opcode_type, 16#09#),
      3215 => to_slv(opcode_type, 16#0F#),
      3216 => to_slv(opcode_type, 16#0E#),
      3217 => to_slv(opcode_type, 16#09#),
      3218 => to_slv(opcode_type, 16#01#),
      3219 => to_slv(opcode_type, 16#0D#),
      3220 => to_slv(opcode_type, 16#0E#),
      3221 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#03#),
      3234 => to_slv(opcode_type, 16#02#),
      3235 => to_slv(opcode_type, 16#09#),
      3236 => to_slv(opcode_type, 16#0E#),
      3237 => to_slv(opcode_type, 16#0B#),
      3238 => to_slv(opcode_type, 16#07#),
      3239 => to_slv(opcode_type, 16#09#),
      3240 => to_slv(opcode_type, 16#07#),
      3241 => to_slv(opcode_type, 16#0A#),
      3242 => to_slv(opcode_type, 16#11#),
      3243 => to_slv(opcode_type, 16#08#),
      3244 => to_slv(opcode_type, 16#0B#),
      3245 => to_slv(opcode_type, 16#0A#),
      3246 => to_slv(opcode_type, 16#06#),
      3247 => to_slv(opcode_type, 16#07#),
      3248 => to_slv(opcode_type, 16#0F#),
      3249 => to_slv(opcode_type, 16#0F#),
      3250 => to_slv(opcode_type, 16#07#),
      3251 => to_slv(opcode_type, 16#0C#),
      3252 => to_slv(opcode_type, 16#0D#),
      3253 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#08#),
      3265 => to_slv(opcode_type, 16#01#),
      3266 => to_slv(opcode_type, 16#07#),
      3267 => to_slv(opcode_type, 16#01#),
      3268 => to_slv(opcode_type, 16#0D#),
      3269 => to_slv(opcode_type, 16#07#),
      3270 => to_slv(opcode_type, 16#0A#),
      3271 => to_slv(opcode_type, 16#0A#),
      3272 => to_slv(opcode_type, 16#06#),
      3273 => to_slv(opcode_type, 16#09#),
      3274 => to_slv(opcode_type, 16#09#),
      3275 => to_slv(opcode_type, 16#D9#),
      3276 => to_slv(opcode_type, 16#10#),
      3277 => to_slv(opcode_type, 16#07#),
      3278 => to_slv(opcode_type, 16#BD#),
      3279 => to_slv(opcode_type, 16#0B#),
      3280 => to_slv(opcode_type, 16#09#),
      3281 => to_slv(opcode_type, 16#08#),
      3282 => to_slv(opcode_type, 16#0B#),
      3283 => to_slv(opcode_type, 16#0F#),
      3284 => to_slv(opcode_type, 16#0F#),
      3285 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#07#),
      3297 => to_slv(opcode_type, 16#03#),
      3298 => to_slv(opcode_type, 16#09#),
      3299 => to_slv(opcode_type, 16#07#),
      3300 => to_slv(opcode_type, 16#31#),
      3301 => to_slv(opcode_type, 16#0D#),
      3302 => to_slv(opcode_type, 16#02#),
      3303 => to_slv(opcode_type, 16#0B#),
      3304 => to_slv(opcode_type, 16#08#),
      3305 => to_slv(opcode_type, 16#08#),
      3306 => to_slv(opcode_type, 16#03#),
      3307 => to_slv(opcode_type, 16#0D#),
      3308 => to_slv(opcode_type, 16#08#),
      3309 => to_slv(opcode_type, 16#0C#),
      3310 => to_slv(opcode_type, 16#0B#),
      3311 => to_slv(opcode_type, 16#08#),
      3312 => to_slv(opcode_type, 16#06#),
      3313 => to_slv(opcode_type, 16#11#),
      3314 => to_slv(opcode_type, 16#0D#),
      3315 => to_slv(opcode_type, 16#04#),
      3316 => to_slv(opcode_type, 16#FC#),
      3317 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#07#),
      3329 => to_slv(opcode_type, 16#03#),
      3330 => to_slv(opcode_type, 16#09#),
      3331 => to_slv(opcode_type, 16#07#),
      3332 => to_slv(opcode_type, 16#10#),
      3333 => to_slv(opcode_type, 16#0F#),
      3334 => to_slv(opcode_type, 16#08#),
      3335 => to_slv(opcode_type, 16#0F#),
      3336 => to_slv(opcode_type, 16#11#),
      3337 => to_slv(opcode_type, 16#08#),
      3338 => to_slv(opcode_type, 16#06#),
      3339 => to_slv(opcode_type, 16#09#),
      3340 => to_slv(opcode_type, 16#10#),
      3341 => to_slv(opcode_type, 16#0B#),
      3342 => to_slv(opcode_type, 16#09#),
      3343 => to_slv(opcode_type, 16#0D#),
      3344 => to_slv(opcode_type, 16#0C#),
      3345 => to_slv(opcode_type, 16#06#),
      3346 => to_slv(opcode_type, 16#02#),
      3347 => to_slv(opcode_type, 16#0E#),
      3348 => to_slv(opcode_type, 16#0D#),
      3349 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#06#),
      3361 => to_slv(opcode_type, 16#06#),
      3362 => to_slv(opcode_type, 16#03#),
      3363 => to_slv(opcode_type, 16#07#),
      3364 => to_slv(opcode_type, 16#9A#),
      3365 => to_slv(opcode_type, 16#0F#),
      3366 => to_slv(opcode_type, 16#04#),
      3367 => to_slv(opcode_type, 16#09#),
      3368 => to_slv(opcode_type, 16#10#),
      3369 => to_slv(opcode_type, 16#0E#),
      3370 => to_slv(opcode_type, 16#09#),
      3371 => to_slv(opcode_type, 16#07#),
      3372 => to_slv(opcode_type, 16#09#),
      3373 => to_slv(opcode_type, 16#0E#),
      3374 => to_slv(opcode_type, 16#E6#),
      3375 => to_slv(opcode_type, 16#09#),
      3376 => to_slv(opcode_type, 16#0D#),
      3377 => to_slv(opcode_type, 16#10#),
      3378 => to_slv(opcode_type, 16#07#),
      3379 => to_slv(opcode_type, 16#10#),
      3380 => to_slv(opcode_type, 16#0A#),
      3381 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#09#),
      3393 => to_slv(opcode_type, 16#08#),
      3394 => to_slv(opcode_type, 16#07#),
      3395 => to_slv(opcode_type, 16#05#),
      3396 => to_slv(opcode_type, 16#10#),
      3397 => to_slv(opcode_type, 16#04#),
      3398 => to_slv(opcode_type, 16#0C#),
      3399 => to_slv(opcode_type, 16#08#),
      3400 => to_slv(opcode_type, 16#03#),
      3401 => to_slv(opcode_type, 16#BC#),
      3402 => to_slv(opcode_type, 16#07#),
      3403 => to_slv(opcode_type, 16#10#),
      3404 => to_slv(opcode_type, 16#0A#),
      3405 => to_slv(opcode_type, 16#06#),
      3406 => to_slv(opcode_type, 16#08#),
      3407 => to_slv(opcode_type, 16#08#),
      3408 => to_slv(opcode_type, 16#0F#),
      3409 => to_slv(opcode_type, 16#0A#),
      3410 => to_slv(opcode_type, 16#05#),
      3411 => to_slv(opcode_type, 16#0B#),
      3412 => to_slv(opcode_type, 16#10#),
      3413 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#04#),
      3426 => to_slv(opcode_type, 16#05#),
      3427 => to_slv(opcode_type, 16#08#),
      3428 => to_slv(opcode_type, 16#0C#),
      3429 => to_slv(opcode_type, 16#0A#),
      3430 => to_slv(opcode_type, 16#08#),
      3431 => to_slv(opcode_type, 16#07#),
      3432 => to_slv(opcode_type, 16#07#),
      3433 => to_slv(opcode_type, 16#33#),
      3434 => to_slv(opcode_type, 16#0F#),
      3435 => to_slv(opcode_type, 16#08#),
      3436 => to_slv(opcode_type, 16#0F#),
      3437 => to_slv(opcode_type, 16#0A#),
      3438 => to_slv(opcode_type, 16#08#),
      3439 => to_slv(opcode_type, 16#08#),
      3440 => to_slv(opcode_type, 16#11#),
      3441 => to_slv(opcode_type, 16#0D#),
      3442 => to_slv(opcode_type, 16#06#),
      3443 => to_slv(opcode_type, 16#0F#),
      3444 => to_slv(opcode_type, 16#11#),
      3445 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#09#),
      3457 => to_slv(opcode_type, 16#09#),
      3458 => to_slv(opcode_type, 16#05#),
      3459 => to_slv(opcode_type, 16#06#),
      3460 => to_slv(opcode_type, 16#0D#),
      3461 => to_slv(opcode_type, 16#0E#),
      3462 => to_slv(opcode_type, 16#04#),
      3463 => to_slv(opcode_type, 16#06#),
      3464 => to_slv(opcode_type, 16#0F#),
      3465 => to_slv(opcode_type, 16#10#),
      3466 => to_slv(opcode_type, 16#09#),
      3467 => to_slv(opcode_type, 16#07#),
      3468 => to_slv(opcode_type, 16#07#),
      3469 => to_slv(opcode_type, 16#10#),
      3470 => to_slv(opcode_type, 16#0B#),
      3471 => to_slv(opcode_type, 16#05#),
      3472 => to_slv(opcode_type, 16#0C#),
      3473 => to_slv(opcode_type, 16#01#),
      3474 => to_slv(opcode_type, 16#07#),
      3475 => to_slv(opcode_type, 16#0E#),
      3476 => to_slv(opcode_type, 16#5A#),
      3477 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#09#),
      3489 => to_slv(opcode_type, 16#01#),
      3490 => to_slv(opcode_type, 16#05#),
      3491 => to_slv(opcode_type, 16#07#),
      3492 => to_slv(opcode_type, 16#0A#),
      3493 => to_slv(opcode_type, 16#76#),
      3494 => to_slv(opcode_type, 16#07#),
      3495 => to_slv(opcode_type, 16#07#),
      3496 => to_slv(opcode_type, 16#09#),
      3497 => to_slv(opcode_type, 16#0D#),
      3498 => to_slv(opcode_type, 16#0A#),
      3499 => to_slv(opcode_type, 16#06#),
      3500 => to_slv(opcode_type, 16#0B#),
      3501 => to_slv(opcode_type, 16#0F#),
      3502 => to_slv(opcode_type, 16#09#),
      3503 => to_slv(opcode_type, 16#08#),
      3504 => to_slv(opcode_type, 16#0E#),
      3505 => to_slv(opcode_type, 16#0C#),
      3506 => to_slv(opcode_type, 16#08#),
      3507 => to_slv(opcode_type, 16#0D#),
      3508 => to_slv(opcode_type, 16#0E#),
      3509 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#09#),
      3521 => to_slv(opcode_type, 16#08#),
      3522 => to_slv(opcode_type, 16#06#),
      3523 => to_slv(opcode_type, 16#02#),
      3524 => to_slv(opcode_type, 16#0F#),
      3525 => to_slv(opcode_type, 16#06#),
      3526 => to_slv(opcode_type, 16#10#),
      3527 => to_slv(opcode_type, 16#0F#),
      3528 => to_slv(opcode_type, 16#03#),
      3529 => to_slv(opcode_type, 16#05#),
      3530 => to_slv(opcode_type, 16#11#),
      3531 => to_slv(opcode_type, 16#08#),
      3532 => to_slv(opcode_type, 16#01#),
      3533 => to_slv(opcode_type, 16#08#),
      3534 => to_slv(opcode_type, 16#0E#),
      3535 => to_slv(opcode_type, 16#10#),
      3536 => to_slv(opcode_type, 16#07#),
      3537 => to_slv(opcode_type, 16#02#),
      3538 => to_slv(opcode_type, 16#0B#),
      3539 => to_slv(opcode_type, 16#03#),
      3540 => to_slv(opcode_type, 16#0E#),
      3541 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#07#),
      3553 => to_slv(opcode_type, 16#04#),
      3554 => to_slv(opcode_type, 16#03#),
      3555 => to_slv(opcode_type, 16#06#),
      3556 => to_slv(opcode_type, 16#11#),
      3557 => to_slv(opcode_type, 16#0F#),
      3558 => to_slv(opcode_type, 16#07#),
      3559 => to_slv(opcode_type, 16#08#),
      3560 => to_slv(opcode_type, 16#06#),
      3561 => to_slv(opcode_type, 16#0C#),
      3562 => to_slv(opcode_type, 16#0E#),
      3563 => to_slv(opcode_type, 16#08#),
      3564 => to_slv(opcode_type, 16#0A#),
      3565 => to_slv(opcode_type, 16#11#),
      3566 => to_slv(opcode_type, 16#06#),
      3567 => to_slv(opcode_type, 16#08#),
      3568 => to_slv(opcode_type, 16#0A#),
      3569 => to_slv(opcode_type, 16#21#),
      3570 => to_slv(opcode_type, 16#07#),
      3571 => to_slv(opcode_type, 16#B7#),
      3572 => to_slv(opcode_type, 16#E7#),
      3573 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#08#),
      3585 => to_slv(opcode_type, 16#09#),
      3586 => to_slv(opcode_type, 16#01#),
      3587 => to_slv(opcode_type, 16#03#),
      3588 => to_slv(opcode_type, 16#10#),
      3589 => to_slv(opcode_type, 16#02#),
      3590 => to_slv(opcode_type, 16#07#),
      3591 => to_slv(opcode_type, 16#10#),
      3592 => to_slv(opcode_type, 16#11#),
      3593 => to_slv(opcode_type, 16#09#),
      3594 => to_slv(opcode_type, 16#09#),
      3595 => to_slv(opcode_type, 16#07#),
      3596 => to_slv(opcode_type, 16#0C#),
      3597 => to_slv(opcode_type, 16#11#),
      3598 => to_slv(opcode_type, 16#01#),
      3599 => to_slv(opcode_type, 16#0B#),
      3600 => to_slv(opcode_type, 16#07#),
      3601 => to_slv(opcode_type, 16#07#),
      3602 => to_slv(opcode_type, 16#0D#),
      3603 => to_slv(opcode_type, 16#0B#),
      3604 => to_slv(opcode_type, 16#0D#),
      3605 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#07#),
      3617 => to_slv(opcode_type, 16#01#),
      3618 => to_slv(opcode_type, 16#05#),
      3619 => to_slv(opcode_type, 16#09#),
      3620 => to_slv(opcode_type, 16#0C#),
      3621 => to_slv(opcode_type, 16#0E#),
      3622 => to_slv(opcode_type, 16#08#),
      3623 => to_slv(opcode_type, 16#07#),
      3624 => to_slv(opcode_type, 16#09#),
      3625 => to_slv(opcode_type, 16#4D#),
      3626 => to_slv(opcode_type, 16#0D#),
      3627 => to_slv(opcode_type, 16#06#),
      3628 => to_slv(opcode_type, 16#0F#),
      3629 => to_slv(opcode_type, 16#0D#),
      3630 => to_slv(opcode_type, 16#08#),
      3631 => to_slv(opcode_type, 16#09#),
      3632 => to_slv(opcode_type, 16#0A#),
      3633 => to_slv(opcode_type, 16#11#),
      3634 => to_slv(opcode_type, 16#08#),
      3635 => to_slv(opcode_type, 16#0F#),
      3636 => to_slv(opcode_type, 16#10#),
      3637 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#07#),
      3649 => to_slv(opcode_type, 16#09#),
      3650 => to_slv(opcode_type, 16#04#),
      3651 => to_slv(opcode_type, 16#04#),
      3652 => to_slv(opcode_type, 16#0A#),
      3653 => to_slv(opcode_type, 16#09#),
      3654 => to_slv(opcode_type, 16#08#),
      3655 => to_slv(opcode_type, 16#0D#),
      3656 => to_slv(opcode_type, 16#10#),
      3657 => to_slv(opcode_type, 16#09#),
      3658 => to_slv(opcode_type, 16#0E#),
      3659 => to_slv(opcode_type, 16#0A#),
      3660 => to_slv(opcode_type, 16#06#),
      3661 => to_slv(opcode_type, 16#03#),
      3662 => to_slv(opcode_type, 16#05#),
      3663 => to_slv(opcode_type, 16#0A#),
      3664 => to_slv(opcode_type, 16#08#),
      3665 => to_slv(opcode_type, 16#06#),
      3666 => to_slv(opcode_type, 16#11#),
      3667 => to_slv(opcode_type, 16#10#),
      3668 => to_slv(opcode_type, 16#0B#),
      3669 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#08#),
      3681 => to_slv(opcode_type, 16#08#),
      3682 => to_slv(opcode_type, 16#03#),
      3683 => to_slv(opcode_type, 16#01#),
      3684 => to_slv(opcode_type, 16#0B#),
      3685 => to_slv(opcode_type, 16#08#),
      3686 => to_slv(opcode_type, 16#09#),
      3687 => to_slv(opcode_type, 16#0F#),
      3688 => to_slv(opcode_type, 16#0C#),
      3689 => to_slv(opcode_type, 16#04#),
      3690 => to_slv(opcode_type, 16#11#),
      3691 => to_slv(opcode_type, 16#07#),
      3692 => to_slv(opcode_type, 16#03#),
      3693 => to_slv(opcode_type, 16#07#),
      3694 => to_slv(opcode_type, 16#0B#),
      3695 => to_slv(opcode_type, 16#0A#),
      3696 => to_slv(opcode_type, 16#06#),
      3697 => to_slv(opcode_type, 16#01#),
      3698 => to_slv(opcode_type, 16#0F#),
      3699 => to_slv(opcode_type, 16#03#),
      3700 => to_slv(opcode_type, 16#0F#),
      3701 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#09#),
      3713 => to_slv(opcode_type, 16#06#),
      3714 => to_slv(opcode_type, 16#05#),
      3715 => to_slv(opcode_type, 16#01#),
      3716 => to_slv(opcode_type, 16#0F#),
      3717 => to_slv(opcode_type, 16#09#),
      3718 => to_slv(opcode_type, 16#01#),
      3719 => to_slv(opcode_type, 16#31#),
      3720 => to_slv(opcode_type, 16#09#),
      3721 => to_slv(opcode_type, 16#10#),
      3722 => to_slv(opcode_type, 16#10#),
      3723 => to_slv(opcode_type, 16#08#),
      3724 => to_slv(opcode_type, 16#04#),
      3725 => to_slv(opcode_type, 16#05#),
      3726 => to_slv(opcode_type, 16#11#),
      3727 => to_slv(opcode_type, 16#08#),
      3728 => to_slv(opcode_type, 16#03#),
      3729 => to_slv(opcode_type, 16#3A#),
      3730 => to_slv(opcode_type, 16#06#),
      3731 => to_slv(opcode_type, 16#11#),
      3732 => to_slv(opcode_type, 16#0D#),
      3733 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#08#),
      3745 => to_slv(opcode_type, 16#07#),
      3746 => to_slv(opcode_type, 16#08#),
      3747 => to_slv(opcode_type, 16#03#),
      3748 => to_slv(opcode_type, 16#11#),
      3749 => to_slv(opcode_type, 16#01#),
      3750 => to_slv(opcode_type, 16#0C#),
      3751 => to_slv(opcode_type, 16#05#),
      3752 => to_slv(opcode_type, 16#05#),
      3753 => to_slv(opcode_type, 16#E6#),
      3754 => to_slv(opcode_type, 16#07#),
      3755 => to_slv(opcode_type, 16#08#),
      3756 => to_slv(opcode_type, 16#04#),
      3757 => to_slv(opcode_type, 16#0B#),
      3758 => to_slv(opcode_type, 16#01#),
      3759 => to_slv(opcode_type, 16#49#),
      3760 => to_slv(opcode_type, 16#07#),
      3761 => to_slv(opcode_type, 16#08#),
      3762 => to_slv(opcode_type, 16#10#),
      3763 => to_slv(opcode_type, 16#0F#),
      3764 => to_slv(opcode_type, 16#E2#),
      3765 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#07#),
      3777 => to_slv(opcode_type, 16#05#),
      3778 => to_slv(opcode_type, 16#04#),
      3779 => to_slv(opcode_type, 16#06#),
      3780 => to_slv(opcode_type, 16#39#),
      3781 => to_slv(opcode_type, 16#10#),
      3782 => to_slv(opcode_type, 16#06#),
      3783 => to_slv(opcode_type, 16#09#),
      3784 => to_slv(opcode_type, 16#06#),
      3785 => to_slv(opcode_type, 16#0B#),
      3786 => to_slv(opcode_type, 16#0D#),
      3787 => to_slv(opcode_type, 16#06#),
      3788 => to_slv(opcode_type, 16#0E#),
      3789 => to_slv(opcode_type, 16#0F#),
      3790 => to_slv(opcode_type, 16#06#),
      3791 => to_slv(opcode_type, 16#08#),
      3792 => to_slv(opcode_type, 16#0A#),
      3793 => to_slv(opcode_type, 16#11#),
      3794 => to_slv(opcode_type, 16#08#),
      3795 => to_slv(opcode_type, 16#0E#),
      3796 => to_slv(opcode_type, 16#0A#),
      3797 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#07#),
      3809 => to_slv(opcode_type, 16#03#),
      3810 => to_slv(opcode_type, 16#05#),
      3811 => to_slv(opcode_type, 16#06#),
      3812 => to_slv(opcode_type, 16#0C#),
      3813 => to_slv(opcode_type, 16#0F#),
      3814 => to_slv(opcode_type, 16#08#),
      3815 => to_slv(opcode_type, 16#09#),
      3816 => to_slv(opcode_type, 16#07#),
      3817 => to_slv(opcode_type, 16#14#),
      3818 => to_slv(opcode_type, 16#0C#),
      3819 => to_slv(opcode_type, 16#09#),
      3820 => to_slv(opcode_type, 16#0B#),
      3821 => to_slv(opcode_type, 16#0F#),
      3822 => to_slv(opcode_type, 16#06#),
      3823 => to_slv(opcode_type, 16#06#),
      3824 => to_slv(opcode_type, 16#0C#),
      3825 => to_slv(opcode_type, 16#0B#),
      3826 => to_slv(opcode_type, 16#07#),
      3827 => to_slv(opcode_type, 16#0D#),
      3828 => to_slv(opcode_type, 16#0E#),
      3829 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#09#),
      3841 => to_slv(opcode_type, 16#06#),
      3842 => to_slv(opcode_type, 16#09#),
      3843 => to_slv(opcode_type, 16#02#),
      3844 => to_slv(opcode_type, 16#0E#),
      3845 => to_slv(opcode_type, 16#06#),
      3846 => to_slv(opcode_type, 16#10#),
      3847 => to_slv(opcode_type, 16#0F#),
      3848 => to_slv(opcode_type, 16#05#),
      3849 => to_slv(opcode_type, 16#06#),
      3850 => to_slv(opcode_type, 16#0B#),
      3851 => to_slv(opcode_type, 16#0D#),
      3852 => to_slv(opcode_type, 16#06#),
      3853 => to_slv(opcode_type, 16#08#),
      3854 => to_slv(opcode_type, 16#09#),
      3855 => to_slv(opcode_type, 16#0D#),
      3856 => to_slv(opcode_type, 16#0D#),
      3857 => to_slv(opcode_type, 16#01#),
      3858 => to_slv(opcode_type, 16#0B#),
      3859 => to_slv(opcode_type, 16#02#),
      3860 => to_slv(opcode_type, 16#10#),
      3861 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#08#),
      3873 => to_slv(opcode_type, 16#06#),
      3874 => to_slv(opcode_type, 16#01#),
      3875 => to_slv(opcode_type, 16#03#),
      3876 => to_slv(opcode_type, 16#0D#),
      3877 => to_slv(opcode_type, 16#04#),
      3878 => to_slv(opcode_type, 16#09#),
      3879 => to_slv(opcode_type, 16#0A#),
      3880 => to_slv(opcode_type, 16#0F#),
      3881 => to_slv(opcode_type, 16#09#),
      3882 => to_slv(opcode_type, 16#03#),
      3883 => to_slv(opcode_type, 16#07#),
      3884 => to_slv(opcode_type, 16#0A#),
      3885 => to_slv(opcode_type, 16#0B#),
      3886 => to_slv(opcode_type, 16#09#),
      3887 => to_slv(opcode_type, 16#07#),
      3888 => to_slv(opcode_type, 16#0B#),
      3889 => to_slv(opcode_type, 16#0C#),
      3890 => to_slv(opcode_type, 16#07#),
      3891 => to_slv(opcode_type, 16#0C#),
      3892 => to_slv(opcode_type, 16#0C#),
      3893 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#07#),
      3905 => to_slv(opcode_type, 16#03#),
      3906 => to_slv(opcode_type, 16#07#),
      3907 => to_slv(opcode_type, 16#02#),
      3908 => to_slv(opcode_type, 16#10#),
      3909 => to_slv(opcode_type, 16#03#),
      3910 => to_slv(opcode_type, 16#0B#),
      3911 => to_slv(opcode_type, 16#09#),
      3912 => to_slv(opcode_type, 16#07#),
      3913 => to_slv(opcode_type, 16#02#),
      3914 => to_slv(opcode_type, 16#EC#),
      3915 => to_slv(opcode_type, 16#08#),
      3916 => to_slv(opcode_type, 16#0E#),
      3917 => to_slv(opcode_type, 16#36#),
      3918 => to_slv(opcode_type, 16#09#),
      3919 => to_slv(opcode_type, 16#07#),
      3920 => to_slv(opcode_type, 16#0F#),
      3921 => to_slv(opcode_type, 16#11#),
      3922 => to_slv(opcode_type, 16#07#),
      3923 => to_slv(opcode_type, 16#11#),
      3924 => to_slv(opcode_type, 16#0C#),
      3925 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#08#),
      3937 => to_slv(opcode_type, 16#02#),
      3938 => to_slv(opcode_type, 16#07#),
      3939 => to_slv(opcode_type, 16#07#),
      3940 => to_slv(opcode_type, 16#10#),
      3941 => to_slv(opcode_type, 16#0B#),
      3942 => to_slv(opcode_type, 16#09#),
      3943 => to_slv(opcode_type, 16#9F#),
      3944 => to_slv(opcode_type, 16#0A#),
      3945 => to_slv(opcode_type, 16#09#),
      3946 => to_slv(opcode_type, 16#09#),
      3947 => to_slv(opcode_type, 16#09#),
      3948 => to_slv(opcode_type, 16#0E#),
      3949 => to_slv(opcode_type, 16#0D#),
      3950 => to_slv(opcode_type, 16#07#),
      3951 => to_slv(opcode_type, 16#10#),
      3952 => to_slv(opcode_type, 16#0F#),
      3953 => to_slv(opcode_type, 16#05#),
      3954 => to_slv(opcode_type, 16#07#),
      3955 => to_slv(opcode_type, 16#0C#),
      3956 => to_slv(opcode_type, 16#0F#),
      3957 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#06#),
      3969 => to_slv(opcode_type, 16#07#),
      3970 => to_slv(opcode_type, 16#09#),
      3971 => to_slv(opcode_type, 16#06#),
      3972 => to_slv(opcode_type, 16#0E#),
      3973 => to_slv(opcode_type, 16#0B#),
      3974 => to_slv(opcode_type, 16#08#),
      3975 => to_slv(opcode_type, 16#0A#),
      3976 => to_slv(opcode_type, 16#7D#),
      3977 => to_slv(opcode_type, 16#05#),
      3978 => to_slv(opcode_type, 16#06#),
      3979 => to_slv(opcode_type, 16#0E#),
      3980 => to_slv(opcode_type, 16#0B#),
      3981 => to_slv(opcode_type, 16#01#),
      3982 => to_slv(opcode_type, 16#08#),
      3983 => to_slv(opcode_type, 16#08#),
      3984 => to_slv(opcode_type, 16#11#),
      3985 => to_slv(opcode_type, 16#0C#),
      3986 => to_slv(opcode_type, 16#07#),
      3987 => to_slv(opcode_type, 16#0F#),
      3988 => to_slv(opcode_type, 16#0D#),
      3989 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#09#),
      4001 => to_slv(opcode_type, 16#02#),
      4002 => to_slv(opcode_type, 16#09#),
      4003 => to_slv(opcode_type, 16#04#),
      4004 => to_slv(opcode_type, 16#0E#),
      4005 => to_slv(opcode_type, 16#02#),
      4006 => to_slv(opcode_type, 16#0E#),
      4007 => to_slv(opcode_type, 16#09#),
      4008 => to_slv(opcode_type, 16#08#),
      4009 => to_slv(opcode_type, 16#07#),
      4010 => to_slv(opcode_type, 16#0B#),
      4011 => to_slv(opcode_type, 16#0F#),
      4012 => to_slv(opcode_type, 16#09#),
      4013 => to_slv(opcode_type, 16#10#),
      4014 => to_slv(opcode_type, 16#4C#),
      4015 => to_slv(opcode_type, 16#09#),
      4016 => to_slv(opcode_type, 16#09#),
      4017 => to_slv(opcode_type, 16#11#),
      4018 => to_slv(opcode_type, 16#0D#),
      4019 => to_slv(opcode_type, 16#03#),
      4020 => to_slv(opcode_type, 16#0D#),
      4021 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#07#),
      4033 => to_slv(opcode_type, 16#07#),
      4034 => to_slv(opcode_type, 16#07#),
      4035 => to_slv(opcode_type, 16#02#),
      4036 => to_slv(opcode_type, 16#0E#),
      4037 => to_slv(opcode_type, 16#05#),
      4038 => to_slv(opcode_type, 16#0A#),
      4039 => to_slv(opcode_type, 16#02#),
      4040 => to_slv(opcode_type, 16#05#),
      4041 => to_slv(opcode_type, 16#0B#),
      4042 => to_slv(opcode_type, 16#08#),
      4043 => to_slv(opcode_type, 16#01#),
      4044 => to_slv(opcode_type, 16#08#),
      4045 => to_slv(opcode_type, 16#0F#),
      4046 => to_slv(opcode_type, 16#85#),
      4047 => to_slv(opcode_type, 16#07#),
      4048 => to_slv(opcode_type, 16#02#),
      4049 => to_slv(opcode_type, 16#11#),
      4050 => to_slv(opcode_type, 16#08#),
      4051 => to_slv(opcode_type, 16#0D#),
      4052 => to_slv(opcode_type, 16#0E#),
      4053 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#04#),
      4066 => to_slv(opcode_type, 16#05#),
      4067 => to_slv(opcode_type, 16#09#),
      4068 => to_slv(opcode_type, 16#0D#),
      4069 => to_slv(opcode_type, 16#0B#),
      4070 => to_slv(opcode_type, 16#06#),
      4071 => to_slv(opcode_type, 16#06#),
      4072 => to_slv(opcode_type, 16#09#),
      4073 => to_slv(opcode_type, 16#0A#),
      4074 => to_slv(opcode_type, 16#0F#),
      4075 => to_slv(opcode_type, 16#07#),
      4076 => to_slv(opcode_type, 16#0F#),
      4077 => to_slv(opcode_type, 16#0E#),
      4078 => to_slv(opcode_type, 16#06#),
      4079 => to_slv(opcode_type, 16#06#),
      4080 => to_slv(opcode_type, 16#11#),
      4081 => to_slv(opcode_type, 16#0C#),
      4082 => to_slv(opcode_type, 16#06#),
      4083 => to_slv(opcode_type, 16#11#),
      4084 => to_slv(opcode_type, 16#0D#),
      4085 to 4095 => (others => '0')
  ),

    -- Bin `22`...
    21 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#08#),
      1 => to_slv(opcode_type, 16#01#),
      2 => to_slv(opcode_type, 16#09#),
      3 => to_slv(opcode_type, 16#06#),
      4 => to_slv(opcode_type, 16#10#),
      5 => to_slv(opcode_type, 16#0D#),
      6 => to_slv(opcode_type, 16#08#),
      7 => to_slv(opcode_type, 16#0C#),
      8 => to_slv(opcode_type, 16#0E#),
      9 => to_slv(opcode_type, 16#08#),
      10 => to_slv(opcode_type, 16#08#),
      11 => to_slv(opcode_type, 16#02#),
      12 => to_slv(opcode_type, 16#0A#),
      13 => to_slv(opcode_type, 16#02#),
      14 => to_slv(opcode_type, 16#0D#),
      15 => to_slv(opcode_type, 16#06#),
      16 => to_slv(opcode_type, 16#07#),
      17 => to_slv(opcode_type, 16#24#),
      18 => to_slv(opcode_type, 16#0A#),
      19 => to_slv(opcode_type, 16#09#),
      20 => to_slv(opcode_type, 16#0C#),
      21 => to_slv(opcode_type, 16#7A#),
      22 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#06#),
      33 => to_slv(opcode_type, 16#05#),
      34 => to_slv(opcode_type, 16#08#),
      35 => to_slv(opcode_type, 16#05#),
      36 => to_slv(opcode_type, 16#11#),
      37 => to_slv(opcode_type, 16#01#),
      38 => to_slv(opcode_type, 16#0E#),
      39 => to_slv(opcode_type, 16#07#),
      40 => to_slv(opcode_type, 16#09#),
      41 => to_slv(opcode_type, 16#07#),
      42 => to_slv(opcode_type, 16#0D#),
      43 => to_slv(opcode_type, 16#24#),
      44 => to_slv(opcode_type, 16#08#),
      45 => to_slv(opcode_type, 16#A1#),
      46 => to_slv(opcode_type, 16#10#),
      47 => to_slv(opcode_type, 16#08#),
      48 => to_slv(opcode_type, 16#07#),
      49 => to_slv(opcode_type, 16#0B#),
      50 => to_slv(opcode_type, 16#CF#),
      51 => to_slv(opcode_type, 16#08#),
      52 => to_slv(opcode_type, 16#0F#),
      53 => to_slv(opcode_type, 16#0C#),
      54 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#08#),
      65 => to_slv(opcode_type, 16#09#),
      66 => to_slv(opcode_type, 16#09#),
      67 => to_slv(opcode_type, 16#06#),
      68 => to_slv(opcode_type, 16#0F#),
      69 => to_slv(opcode_type, 16#0A#),
      70 => to_slv(opcode_type, 16#02#),
      71 => to_slv(opcode_type, 16#0C#),
      72 => to_slv(opcode_type, 16#02#),
      73 => to_slv(opcode_type, 16#04#),
      74 => to_slv(opcode_type, 16#0C#),
      75 => to_slv(opcode_type, 16#09#),
      76 => to_slv(opcode_type, 16#09#),
      77 => to_slv(opcode_type, 16#01#),
      78 => to_slv(opcode_type, 16#0F#),
      79 => to_slv(opcode_type, 16#04#),
      80 => to_slv(opcode_type, 16#0A#),
      81 => to_slv(opcode_type, 16#08#),
      82 => to_slv(opcode_type, 16#08#),
      83 => to_slv(opcode_type, 16#0E#),
      84 => to_slv(opcode_type, 16#0D#),
      85 => to_slv(opcode_type, 16#F6#),
      86 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#09#),
      97 => to_slv(opcode_type, 16#01#),
      98 => to_slv(opcode_type, 16#09#),
      99 => to_slv(opcode_type, 16#03#),
      100 => to_slv(opcode_type, 16#0A#),
      101 => to_slv(opcode_type, 16#09#),
      102 => to_slv(opcode_type, 16#10#),
      103 => to_slv(opcode_type, 16#10#),
      104 => to_slv(opcode_type, 16#07#),
      105 => to_slv(opcode_type, 16#06#),
      106 => to_slv(opcode_type, 16#03#),
      107 => to_slv(opcode_type, 16#0F#),
      108 => to_slv(opcode_type, 16#06#),
      109 => to_slv(opcode_type, 16#0B#),
      110 => to_slv(opcode_type, 16#11#),
      111 => to_slv(opcode_type, 16#06#),
      112 => to_slv(opcode_type, 16#06#),
      113 => to_slv(opcode_type, 16#0D#),
      114 => to_slv(opcode_type, 16#11#),
      115 => to_slv(opcode_type, 16#08#),
      116 => to_slv(opcode_type, 16#0E#),
      117 => to_slv(opcode_type, 16#11#),
      118 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#07#),
      129 => to_slv(opcode_type, 16#08#),
      130 => to_slv(opcode_type, 16#04#),
      131 => to_slv(opcode_type, 16#09#),
      132 => to_slv(opcode_type, 16#0E#),
      133 => to_slv(opcode_type, 16#0B#),
      134 => to_slv(opcode_type, 16#08#),
      135 => to_slv(opcode_type, 16#03#),
      136 => to_slv(opcode_type, 16#0E#),
      137 => to_slv(opcode_type, 16#01#),
      138 => to_slv(opcode_type, 16#0B#),
      139 => to_slv(opcode_type, 16#07#),
      140 => to_slv(opcode_type, 16#07#),
      141 => to_slv(opcode_type, 16#07#),
      142 => to_slv(opcode_type, 16#0A#),
      143 => to_slv(opcode_type, 16#0B#),
      144 => to_slv(opcode_type, 16#07#),
      145 => to_slv(opcode_type, 16#11#),
      146 => to_slv(opcode_type, 16#85#),
      147 => to_slv(opcode_type, 16#09#),
      148 => to_slv(opcode_type, 16#0F#),
      149 => to_slv(opcode_type, 16#0E#),
      150 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#06#),
      161 => to_slv(opcode_type, 16#02#),
      162 => to_slv(opcode_type, 16#09#),
      163 => to_slv(opcode_type, 16#08#),
      164 => to_slv(opcode_type, 16#0F#),
      165 => to_slv(opcode_type, 16#0B#),
      166 => to_slv(opcode_type, 16#05#),
      167 => to_slv(opcode_type, 16#0F#),
      168 => to_slv(opcode_type, 16#09#),
      169 => to_slv(opcode_type, 16#06#),
      170 => to_slv(opcode_type, 16#07#),
      171 => to_slv(opcode_type, 16#0E#),
      172 => to_slv(opcode_type, 16#0A#),
      173 => to_slv(opcode_type, 16#03#),
      174 => to_slv(opcode_type, 16#0C#),
      175 => to_slv(opcode_type, 16#08#),
      176 => to_slv(opcode_type, 16#08#),
      177 => to_slv(opcode_type, 16#0A#),
      178 => to_slv(opcode_type, 16#0D#),
      179 => to_slv(opcode_type, 16#08#),
      180 => to_slv(opcode_type, 16#0D#),
      181 => to_slv(opcode_type, 16#0A#),
      182 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#06#),
      193 => to_slv(opcode_type, 16#07#),
      194 => to_slv(opcode_type, 16#02#),
      195 => to_slv(opcode_type, 16#06#),
      196 => to_slv(opcode_type, 16#10#),
      197 => to_slv(opcode_type, 16#3D#),
      198 => to_slv(opcode_type, 16#07#),
      199 => to_slv(opcode_type, 16#08#),
      200 => to_slv(opcode_type, 16#0E#),
      201 => to_slv(opcode_type, 16#0C#),
      202 => to_slv(opcode_type, 16#01#),
      203 => to_slv(opcode_type, 16#0E#),
      204 => to_slv(opcode_type, 16#07#),
      205 => to_slv(opcode_type, 16#06#),
      206 => to_slv(opcode_type, 16#03#),
      207 => to_slv(opcode_type, 16#0E#),
      208 => to_slv(opcode_type, 16#01#),
      209 => to_slv(opcode_type, 16#0D#),
      210 => to_slv(opcode_type, 16#03#),
      211 => to_slv(opcode_type, 16#08#),
      212 => to_slv(opcode_type, 16#0A#),
      213 => to_slv(opcode_type, 16#11#),
      214 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#07#),
      225 => to_slv(opcode_type, 16#06#),
      226 => to_slv(opcode_type, 16#06#),
      227 => to_slv(opcode_type, 16#07#),
      228 => to_slv(opcode_type, 16#0D#),
      229 => to_slv(opcode_type, 16#A6#),
      230 => to_slv(opcode_type, 16#06#),
      231 => to_slv(opcode_type, 16#0C#),
      232 => to_slv(opcode_type, 16#0E#),
      233 => to_slv(opcode_type, 16#05#),
      234 => to_slv(opcode_type, 16#04#),
      235 => to_slv(opcode_type, 16#0A#),
      236 => to_slv(opcode_type, 16#09#),
      237 => to_slv(opcode_type, 16#04#),
      238 => to_slv(opcode_type, 16#04#),
      239 => to_slv(opcode_type, 16#0B#),
      240 => to_slv(opcode_type, 16#06#),
      241 => to_slv(opcode_type, 16#07#),
      242 => to_slv(opcode_type, 16#0B#),
      243 => to_slv(opcode_type, 16#10#),
      244 => to_slv(opcode_type, 16#05#),
      245 => to_slv(opcode_type, 16#0D#),
      246 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#09#),
      257 => to_slv(opcode_type, 16#04#),
      258 => to_slv(opcode_type, 16#08#),
      259 => to_slv(opcode_type, 16#03#),
      260 => to_slv(opcode_type, 16#0A#),
      261 => to_slv(opcode_type, 16#06#),
      262 => to_slv(opcode_type, 16#0D#),
      263 => to_slv(opcode_type, 16#10#),
      264 => to_slv(opcode_type, 16#09#),
      265 => to_slv(opcode_type, 16#06#),
      266 => to_slv(opcode_type, 16#06#),
      267 => to_slv(opcode_type, 16#D5#),
      268 => to_slv(opcode_type, 16#11#),
      269 => to_slv(opcode_type, 16#09#),
      270 => to_slv(opcode_type, 16#0B#),
      271 => to_slv(opcode_type, 16#0E#),
      272 => to_slv(opcode_type, 16#06#),
      273 => to_slv(opcode_type, 16#09#),
      274 => to_slv(opcode_type, 16#10#),
      275 => to_slv(opcode_type, 16#11#),
      276 => to_slv(opcode_type, 16#03#),
      277 => to_slv(opcode_type, 16#11#),
      278 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#08#),
      289 => to_slv(opcode_type, 16#09#),
      290 => to_slv(opcode_type, 16#04#),
      291 => to_slv(opcode_type, 16#01#),
      292 => to_slv(opcode_type, 16#10#),
      293 => to_slv(opcode_type, 16#07#),
      294 => to_slv(opcode_type, 16#05#),
      295 => to_slv(opcode_type, 16#0F#),
      296 => to_slv(opcode_type, 16#07#),
      297 => to_slv(opcode_type, 16#0A#),
      298 => to_slv(opcode_type, 16#0C#),
      299 => to_slv(opcode_type, 16#09#),
      300 => to_slv(opcode_type, 16#05#),
      301 => to_slv(opcode_type, 16#07#),
      302 => to_slv(opcode_type, 16#0A#),
      303 => to_slv(opcode_type, 16#0D#),
      304 => to_slv(opcode_type, 16#07#),
      305 => to_slv(opcode_type, 16#08#),
      306 => to_slv(opcode_type, 16#10#),
      307 => to_slv(opcode_type, 16#10#),
      308 => to_slv(opcode_type, 16#01#),
      309 => to_slv(opcode_type, 16#0F#),
      310 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#08#),
      321 => to_slv(opcode_type, 16#04#),
      322 => to_slv(opcode_type, 16#08#),
      323 => to_slv(opcode_type, 16#09#),
      324 => to_slv(opcode_type, 16#0D#),
      325 => to_slv(opcode_type, 16#11#),
      326 => to_slv(opcode_type, 16#06#),
      327 => to_slv(opcode_type, 16#0B#),
      328 => to_slv(opcode_type, 16#11#),
      329 => to_slv(opcode_type, 16#06#),
      330 => to_slv(opcode_type, 16#07#),
      331 => to_slv(opcode_type, 16#06#),
      332 => to_slv(opcode_type, 16#0B#),
      333 => to_slv(opcode_type, 16#10#),
      334 => to_slv(opcode_type, 16#05#),
      335 => to_slv(opcode_type, 16#19#),
      336 => to_slv(opcode_type, 16#06#),
      337 => to_slv(opcode_type, 16#01#),
      338 => to_slv(opcode_type, 16#0B#),
      339 => to_slv(opcode_type, 16#07#),
      340 => to_slv(opcode_type, 16#0D#),
      341 => to_slv(opcode_type, 16#0F#),
      342 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#06#),
      353 => to_slv(opcode_type, 16#08#),
      354 => to_slv(opcode_type, 16#04#),
      355 => to_slv(opcode_type, 16#04#),
      356 => to_slv(opcode_type, 16#0A#),
      357 => to_slv(opcode_type, 16#03#),
      358 => to_slv(opcode_type, 16#08#),
      359 => to_slv(opcode_type, 16#0F#),
      360 => to_slv(opcode_type, 16#0F#),
      361 => to_slv(opcode_type, 16#07#),
      362 => to_slv(opcode_type, 16#06#),
      363 => to_slv(opcode_type, 16#05#),
      364 => to_slv(opcode_type, 16#0C#),
      365 => to_slv(opcode_type, 16#03#),
      366 => to_slv(opcode_type, 16#0A#),
      367 => to_slv(opcode_type, 16#09#),
      368 => to_slv(opcode_type, 16#07#),
      369 => to_slv(opcode_type, 16#0D#),
      370 => to_slv(opcode_type, 16#0D#),
      371 => to_slv(opcode_type, 16#06#),
      372 => to_slv(opcode_type, 16#0D#),
      373 => to_slv(opcode_type, 16#0F#),
      374 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#08#),
      385 => to_slv(opcode_type, 16#04#),
      386 => to_slv(opcode_type, 16#06#),
      387 => to_slv(opcode_type, 16#05#),
      388 => to_slv(opcode_type, 16#FF#),
      389 => to_slv(opcode_type, 16#02#),
      390 => to_slv(opcode_type, 16#0E#),
      391 => to_slv(opcode_type, 16#08#),
      392 => to_slv(opcode_type, 16#06#),
      393 => to_slv(opcode_type, 16#08#),
      394 => to_slv(opcode_type, 16#0F#),
      395 => to_slv(opcode_type, 16#0D#),
      396 => to_slv(opcode_type, 16#06#),
      397 => to_slv(opcode_type, 16#0D#),
      398 => to_slv(opcode_type, 16#0B#),
      399 => to_slv(opcode_type, 16#08#),
      400 => to_slv(opcode_type, 16#07#),
      401 => to_slv(opcode_type, 16#11#),
      402 => to_slv(opcode_type, 16#0F#),
      403 => to_slv(opcode_type, 16#08#),
      404 => to_slv(opcode_type, 16#0A#),
      405 => to_slv(opcode_type, 16#0E#),
      406 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#06#),
      417 => to_slv(opcode_type, 16#05#),
      418 => to_slv(opcode_type, 16#08#),
      419 => to_slv(opcode_type, 16#04#),
      420 => to_slv(opcode_type, 16#0A#),
      421 => to_slv(opcode_type, 16#03#),
      422 => to_slv(opcode_type, 16#0E#),
      423 => to_slv(opcode_type, 16#06#),
      424 => to_slv(opcode_type, 16#08#),
      425 => to_slv(opcode_type, 16#08#),
      426 => to_slv(opcode_type, 16#AB#),
      427 => to_slv(opcode_type, 16#10#),
      428 => to_slv(opcode_type, 16#08#),
      429 => to_slv(opcode_type, 16#11#),
      430 => to_slv(opcode_type, 16#0F#),
      431 => to_slv(opcode_type, 16#07#),
      432 => to_slv(opcode_type, 16#08#),
      433 => to_slv(opcode_type, 16#0B#),
      434 => to_slv(opcode_type, 16#0A#),
      435 => to_slv(opcode_type, 16#06#),
      436 => to_slv(opcode_type, 16#0D#),
      437 => to_slv(opcode_type, 16#11#),
      438 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#07#),
      449 => to_slv(opcode_type, 16#03#),
      450 => to_slv(opcode_type, 16#09#),
      451 => to_slv(opcode_type, 16#04#),
      452 => to_slv(opcode_type, 16#0B#),
      453 => to_slv(opcode_type, 16#02#),
      454 => to_slv(opcode_type, 16#BF#),
      455 => to_slv(opcode_type, 16#09#),
      456 => to_slv(opcode_type, 16#08#),
      457 => to_slv(opcode_type, 16#06#),
      458 => to_slv(opcode_type, 16#10#),
      459 => to_slv(opcode_type, 16#10#),
      460 => to_slv(opcode_type, 16#07#),
      461 => to_slv(opcode_type, 16#0B#),
      462 => to_slv(opcode_type, 16#97#),
      463 => to_slv(opcode_type, 16#06#),
      464 => to_slv(opcode_type, 16#07#),
      465 => to_slv(opcode_type, 16#E6#),
      466 => to_slv(opcode_type, 16#0D#),
      467 => to_slv(opcode_type, 16#09#),
      468 => to_slv(opcode_type, 16#0D#),
      469 => to_slv(opcode_type, 16#0B#),
      470 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#06#),
      481 => to_slv(opcode_type, 16#06#),
      482 => to_slv(opcode_type, 16#05#),
      483 => to_slv(opcode_type, 16#01#),
      484 => to_slv(opcode_type, 16#0F#),
      485 => to_slv(opcode_type, 16#05#),
      486 => to_slv(opcode_type, 16#04#),
      487 => to_slv(opcode_type, 16#11#),
      488 => to_slv(opcode_type, 16#07#),
      489 => to_slv(opcode_type, 16#09#),
      490 => to_slv(opcode_type, 16#04#),
      491 => to_slv(opcode_type, 16#10#),
      492 => to_slv(opcode_type, 16#06#),
      493 => to_slv(opcode_type, 16#D3#),
      494 => to_slv(opcode_type, 16#0D#),
      495 => to_slv(opcode_type, 16#07#),
      496 => to_slv(opcode_type, 16#07#),
      497 => to_slv(opcode_type, 16#0F#),
      498 => to_slv(opcode_type, 16#11#),
      499 => to_slv(opcode_type, 16#07#),
      500 => to_slv(opcode_type, 16#0C#),
      501 => to_slv(opcode_type, 16#0F#),
      502 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#04#),
      514 => to_slv(opcode_type, 16#08#),
      515 => to_slv(opcode_type, 16#07#),
      516 => to_slv(opcode_type, 16#10#),
      517 => to_slv(opcode_type, 16#0E#),
      518 => to_slv(opcode_type, 16#02#),
      519 => to_slv(opcode_type, 16#0E#),
      520 => to_slv(opcode_type, 16#09#),
      521 => to_slv(opcode_type, 16#08#),
      522 => to_slv(opcode_type, 16#09#),
      523 => to_slv(opcode_type, 16#10#),
      524 => to_slv(opcode_type, 16#11#),
      525 => to_slv(opcode_type, 16#08#),
      526 => to_slv(opcode_type, 16#42#),
      527 => to_slv(opcode_type, 16#0B#),
      528 => to_slv(opcode_type, 16#08#),
      529 => to_slv(opcode_type, 16#02#),
      530 => to_slv(opcode_type, 16#0E#),
      531 => to_slv(opcode_type, 16#09#),
      532 => to_slv(opcode_type, 16#0F#),
      533 => to_slv(opcode_type, 16#0B#),
      534 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#09#),
      545 => to_slv(opcode_type, 16#08#),
      546 => to_slv(opcode_type, 16#03#),
      547 => to_slv(opcode_type, 16#02#),
      548 => to_slv(opcode_type, 16#0E#),
      549 => to_slv(opcode_type, 16#08#),
      550 => to_slv(opcode_type, 16#08#),
      551 => to_slv(opcode_type, 16#0A#),
      552 => to_slv(opcode_type, 16#10#),
      553 => to_slv(opcode_type, 16#04#),
      554 => to_slv(opcode_type, 16#0E#),
      555 => to_slv(opcode_type, 16#08#),
      556 => to_slv(opcode_type, 16#07#),
      557 => to_slv(opcode_type, 16#04#),
      558 => to_slv(opcode_type, 16#0B#),
      559 => to_slv(opcode_type, 16#07#),
      560 => to_slv(opcode_type, 16#0F#),
      561 => to_slv(opcode_type, 16#11#),
      562 => to_slv(opcode_type, 16#07#),
      563 => to_slv(opcode_type, 16#03#),
      564 => to_slv(opcode_type, 16#11#),
      565 => to_slv(opcode_type, 16#0F#),
      566 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#07#),
      577 => to_slv(opcode_type, 16#02#),
      578 => to_slv(opcode_type, 16#06#),
      579 => to_slv(opcode_type, 16#07#),
      580 => to_slv(opcode_type, 16#DC#),
      581 => to_slv(opcode_type, 16#0F#),
      582 => to_slv(opcode_type, 16#06#),
      583 => to_slv(opcode_type, 16#11#),
      584 => to_slv(opcode_type, 16#10#),
      585 => to_slv(opcode_type, 16#09#),
      586 => to_slv(opcode_type, 16#06#),
      587 => to_slv(opcode_type, 16#07#),
      588 => to_slv(opcode_type, 16#10#),
      589 => to_slv(opcode_type, 16#0D#),
      590 => to_slv(opcode_type, 16#03#),
      591 => to_slv(opcode_type, 16#D6#),
      592 => to_slv(opcode_type, 16#06#),
      593 => to_slv(opcode_type, 16#03#),
      594 => to_slv(opcode_type, 16#0D#),
      595 => to_slv(opcode_type, 16#07#),
      596 => to_slv(opcode_type, 16#0D#),
      597 => to_slv(opcode_type, 16#B1#),
      598 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#06#),
      609 => to_slv(opcode_type, 16#03#),
      610 => to_slv(opcode_type, 16#06#),
      611 => to_slv(opcode_type, 16#05#),
      612 => to_slv(opcode_type, 16#0E#),
      613 => to_slv(opcode_type, 16#02#),
      614 => to_slv(opcode_type, 16#11#),
      615 => to_slv(opcode_type, 16#06#),
      616 => to_slv(opcode_type, 16#06#),
      617 => to_slv(opcode_type, 16#06#),
      618 => to_slv(opcode_type, 16#EE#),
      619 => to_slv(opcode_type, 16#0A#),
      620 => to_slv(opcode_type, 16#08#),
      621 => to_slv(opcode_type, 16#10#),
      622 => to_slv(opcode_type, 16#0E#),
      623 => to_slv(opcode_type, 16#07#),
      624 => to_slv(opcode_type, 16#06#),
      625 => to_slv(opcode_type, 16#10#),
      626 => to_slv(opcode_type, 16#0E#),
      627 => to_slv(opcode_type, 16#08#),
      628 => to_slv(opcode_type, 16#C8#),
      629 => to_slv(opcode_type, 16#0B#),
      630 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#08#),
      641 => to_slv(opcode_type, 16#07#),
      642 => to_slv(opcode_type, 16#06#),
      643 => to_slv(opcode_type, 16#05#),
      644 => to_slv(opcode_type, 16#0A#),
      645 => to_slv(opcode_type, 16#06#),
      646 => to_slv(opcode_type, 16#10#),
      647 => to_slv(opcode_type, 16#10#),
      648 => to_slv(opcode_type, 16#06#),
      649 => to_slv(opcode_type, 16#03#),
      650 => to_slv(opcode_type, 16#0A#),
      651 => to_slv(opcode_type, 16#04#),
      652 => to_slv(opcode_type, 16#CB#),
      653 => to_slv(opcode_type, 16#09#),
      654 => to_slv(opcode_type, 16#07#),
      655 => to_slv(opcode_type, 16#03#),
      656 => to_slv(opcode_type, 16#0E#),
      657 => to_slv(opcode_type, 16#05#),
      658 => to_slv(opcode_type, 16#0B#),
      659 => to_slv(opcode_type, 16#02#),
      660 => to_slv(opcode_type, 16#04#),
      661 => to_slv(opcode_type, 16#10#),
      662 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#09#),
      673 => to_slv(opcode_type, 16#02#),
      674 => to_slv(opcode_type, 16#07#),
      675 => to_slv(opcode_type, 16#09#),
      676 => to_slv(opcode_type, 16#11#),
      677 => to_slv(opcode_type, 16#0D#),
      678 => to_slv(opcode_type, 16#05#),
      679 => to_slv(opcode_type, 16#11#),
      680 => to_slv(opcode_type, 16#07#),
      681 => to_slv(opcode_type, 16#07#),
      682 => to_slv(opcode_type, 16#08#),
      683 => to_slv(opcode_type, 16#11#),
      684 => to_slv(opcode_type, 16#0E#),
      685 => to_slv(opcode_type, 16#09#),
      686 => to_slv(opcode_type, 16#0A#),
      687 => to_slv(opcode_type, 16#0E#),
      688 => to_slv(opcode_type, 16#06#),
      689 => to_slv(opcode_type, 16#01#),
      690 => to_slv(opcode_type, 16#0E#),
      691 => to_slv(opcode_type, 16#09#),
      692 => to_slv(opcode_type, 16#0F#),
      693 => to_slv(opcode_type, 16#0B#),
      694 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#08#),
      705 => to_slv(opcode_type, 16#04#),
      706 => to_slv(opcode_type, 16#08#),
      707 => to_slv(opcode_type, 16#08#),
      708 => to_slv(opcode_type, 16#AF#),
      709 => to_slv(opcode_type, 16#11#),
      710 => to_slv(opcode_type, 16#09#),
      711 => to_slv(opcode_type, 16#0D#),
      712 => to_slv(opcode_type, 16#0A#),
      713 => to_slv(opcode_type, 16#08#),
      714 => to_slv(opcode_type, 16#06#),
      715 => to_slv(opcode_type, 16#03#),
      716 => to_slv(opcode_type, 16#0D#),
      717 => to_slv(opcode_type, 16#03#),
      718 => to_slv(opcode_type, 16#0B#),
      719 => to_slv(opcode_type, 16#09#),
      720 => to_slv(opcode_type, 16#07#),
      721 => to_slv(opcode_type, 16#0D#),
      722 => to_slv(opcode_type, 16#0D#),
      723 => to_slv(opcode_type, 16#09#),
      724 => to_slv(opcode_type, 16#0C#),
      725 => to_slv(opcode_type, 16#0D#),
      726 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#07#),
      737 => to_slv(opcode_type, 16#06#),
      738 => to_slv(opcode_type, 16#09#),
      739 => to_slv(opcode_type, 16#01#),
      740 => to_slv(opcode_type, 16#97#),
      741 => to_slv(opcode_type, 16#03#),
      742 => to_slv(opcode_type, 16#0C#),
      743 => to_slv(opcode_type, 16#01#),
      744 => to_slv(opcode_type, 16#02#),
      745 => to_slv(opcode_type, 16#0D#),
      746 => to_slv(opcode_type, 16#08#),
      747 => to_slv(opcode_type, 16#04#),
      748 => to_slv(opcode_type, 16#07#),
      749 => to_slv(opcode_type, 16#0B#),
      750 => to_slv(opcode_type, 16#11#),
      751 => to_slv(opcode_type, 16#08#),
      752 => to_slv(opcode_type, 16#06#),
      753 => to_slv(opcode_type, 16#0E#),
      754 => to_slv(opcode_type, 16#4E#),
      755 => to_slv(opcode_type, 16#06#),
      756 => to_slv(opcode_type, 16#0A#),
      757 => to_slv(opcode_type, 16#87#),
      758 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#09#),
      769 => to_slv(opcode_type, 16#07#),
      770 => to_slv(opcode_type, 16#02#),
      771 => to_slv(opcode_type, 16#05#),
      772 => to_slv(opcode_type, 16#34#),
      773 => to_slv(opcode_type, 16#05#),
      774 => to_slv(opcode_type, 16#09#),
      775 => to_slv(opcode_type, 16#0A#),
      776 => to_slv(opcode_type, 16#0F#),
      777 => to_slv(opcode_type, 16#07#),
      778 => to_slv(opcode_type, 16#08#),
      779 => to_slv(opcode_type, 16#02#),
      780 => to_slv(opcode_type, 16#0E#),
      781 => to_slv(opcode_type, 16#02#),
      782 => to_slv(opcode_type, 16#0E#),
      783 => to_slv(opcode_type, 16#08#),
      784 => to_slv(opcode_type, 16#08#),
      785 => to_slv(opcode_type, 16#11#),
      786 => to_slv(opcode_type, 16#0E#),
      787 => to_slv(opcode_type, 16#09#),
      788 => to_slv(opcode_type, 16#0A#),
      789 => to_slv(opcode_type, 16#0C#),
      790 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#08#),
      801 => to_slv(opcode_type, 16#09#),
      802 => to_slv(opcode_type, 16#01#),
      803 => to_slv(opcode_type, 16#08#),
      804 => to_slv(opcode_type, 16#0C#),
      805 => to_slv(opcode_type, 16#11#),
      806 => to_slv(opcode_type, 16#04#),
      807 => to_slv(opcode_type, 16#01#),
      808 => to_slv(opcode_type, 16#0B#),
      809 => to_slv(opcode_type, 16#09#),
      810 => to_slv(opcode_type, 16#09#),
      811 => to_slv(opcode_type, 16#03#),
      812 => to_slv(opcode_type, 16#0F#),
      813 => to_slv(opcode_type, 16#03#),
      814 => to_slv(opcode_type, 16#0A#),
      815 => to_slv(opcode_type, 16#09#),
      816 => to_slv(opcode_type, 16#09#),
      817 => to_slv(opcode_type, 16#0D#),
      818 => to_slv(opcode_type, 16#0D#),
      819 => to_slv(opcode_type, 16#06#),
      820 => to_slv(opcode_type, 16#0E#),
      821 => to_slv(opcode_type, 16#10#),
      822 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#07#),
      833 => to_slv(opcode_type, 16#07#),
      834 => to_slv(opcode_type, 16#02#),
      835 => to_slv(opcode_type, 16#08#),
      836 => to_slv(opcode_type, 16#0C#),
      837 => to_slv(opcode_type, 16#11#),
      838 => to_slv(opcode_type, 16#03#),
      839 => to_slv(opcode_type, 16#08#),
      840 => to_slv(opcode_type, 16#0C#),
      841 => to_slv(opcode_type, 16#10#),
      842 => to_slv(opcode_type, 16#09#),
      843 => to_slv(opcode_type, 16#03#),
      844 => to_slv(opcode_type, 16#06#),
      845 => to_slv(opcode_type, 16#0B#),
      846 => to_slv(opcode_type, 16#10#),
      847 => to_slv(opcode_type, 16#07#),
      848 => to_slv(opcode_type, 16#08#),
      849 => to_slv(opcode_type, 16#11#),
      850 => to_slv(opcode_type, 16#0D#),
      851 => to_slv(opcode_type, 16#08#),
      852 => to_slv(opcode_type, 16#A5#),
      853 => to_slv(opcode_type, 16#0B#),
      854 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#06#),
      865 => to_slv(opcode_type, 16#06#),
      866 => to_slv(opcode_type, 16#03#),
      867 => to_slv(opcode_type, 16#05#),
      868 => to_slv(opcode_type, 16#0A#),
      869 => to_slv(opcode_type, 16#06#),
      870 => to_slv(opcode_type, 16#01#),
      871 => to_slv(opcode_type, 16#0E#),
      872 => to_slv(opcode_type, 16#07#),
      873 => to_slv(opcode_type, 16#44#),
      874 => to_slv(opcode_type, 16#11#),
      875 => to_slv(opcode_type, 16#08#),
      876 => to_slv(opcode_type, 16#05#),
      877 => to_slv(opcode_type, 16#06#),
      878 => to_slv(opcode_type, 16#0C#),
      879 => to_slv(opcode_type, 16#0E#),
      880 => to_slv(opcode_type, 16#09#),
      881 => to_slv(opcode_type, 16#01#),
      882 => to_slv(opcode_type, 16#0F#),
      883 => to_slv(opcode_type, 16#06#),
      884 => to_slv(opcode_type, 16#0F#),
      885 => to_slv(opcode_type, 16#0A#),
      886 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#01#),
      898 => to_slv(opcode_type, 16#08#),
      899 => to_slv(opcode_type, 16#03#),
      900 => to_slv(opcode_type, 16#CD#),
      901 => to_slv(opcode_type, 16#07#),
      902 => to_slv(opcode_type, 16#10#),
      903 => to_slv(opcode_type, 16#ED#),
      904 => to_slv(opcode_type, 16#09#),
      905 => to_slv(opcode_type, 16#09#),
      906 => to_slv(opcode_type, 16#01#),
      907 => to_slv(opcode_type, 16#0C#),
      908 => to_slv(opcode_type, 16#07#),
      909 => to_slv(opcode_type, 16#0F#),
      910 => to_slv(opcode_type, 16#10#),
      911 => to_slv(opcode_type, 16#07#),
      912 => to_slv(opcode_type, 16#08#),
      913 => to_slv(opcode_type, 16#0F#),
      914 => to_slv(opcode_type, 16#0F#),
      915 => to_slv(opcode_type, 16#09#),
      916 => to_slv(opcode_type, 16#0A#),
      917 => to_slv(opcode_type, 16#0D#),
      918 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#07#),
      929 => to_slv(opcode_type, 16#06#),
      930 => to_slv(opcode_type, 16#06#),
      931 => to_slv(opcode_type, 16#09#),
      932 => to_slv(opcode_type, 16#DB#),
      933 => to_slv(opcode_type, 16#0B#),
      934 => to_slv(opcode_type, 16#02#),
      935 => to_slv(opcode_type, 16#0C#),
      936 => to_slv(opcode_type, 16#02#),
      937 => to_slv(opcode_type, 16#01#),
      938 => to_slv(opcode_type, 16#0E#),
      939 => to_slv(opcode_type, 16#07#),
      940 => to_slv(opcode_type, 16#04#),
      941 => to_slv(opcode_type, 16#04#),
      942 => to_slv(opcode_type, 16#0D#),
      943 => to_slv(opcode_type, 16#07#),
      944 => to_slv(opcode_type, 16#06#),
      945 => to_slv(opcode_type, 16#10#),
      946 => to_slv(opcode_type, 16#0B#),
      947 => to_slv(opcode_type, 16#08#),
      948 => to_slv(opcode_type, 16#11#),
      949 => to_slv(opcode_type, 16#0C#),
      950 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#06#),
      961 => to_slv(opcode_type, 16#07#),
      962 => to_slv(opcode_type, 16#05#),
      963 => to_slv(opcode_type, 16#08#),
      964 => to_slv(opcode_type, 16#10#),
      965 => to_slv(opcode_type, 16#11#),
      966 => to_slv(opcode_type, 16#07#),
      967 => to_slv(opcode_type, 16#07#),
      968 => to_slv(opcode_type, 16#0C#),
      969 => to_slv(opcode_type, 16#0F#),
      970 => to_slv(opcode_type, 16#01#),
      971 => to_slv(opcode_type, 16#0A#),
      972 => to_slv(opcode_type, 16#07#),
      973 => to_slv(opcode_type, 16#04#),
      974 => to_slv(opcode_type, 16#01#),
      975 => to_slv(opcode_type, 16#11#),
      976 => to_slv(opcode_type, 16#09#),
      977 => to_slv(opcode_type, 16#08#),
      978 => to_slv(opcode_type, 16#0C#),
      979 => to_slv(opcode_type, 16#11#),
      980 => to_slv(opcode_type, 16#05#),
      981 => to_slv(opcode_type, 16#11#),
      982 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#07#),
      993 => to_slv(opcode_type, 16#04#),
      994 => to_slv(opcode_type, 16#08#),
      995 => to_slv(opcode_type, 16#06#),
      996 => to_slv(opcode_type, 16#0A#),
      997 => to_slv(opcode_type, 16#0A#),
      998 => to_slv(opcode_type, 16#01#),
      999 => to_slv(opcode_type, 16#11#),
      1000 => to_slv(opcode_type, 16#06#),
      1001 => to_slv(opcode_type, 16#07#),
      1002 => to_slv(opcode_type, 16#03#),
      1003 => to_slv(opcode_type, 16#11#),
      1004 => to_slv(opcode_type, 16#06#),
      1005 => to_slv(opcode_type, 16#0A#),
      1006 => to_slv(opcode_type, 16#0A#),
      1007 => to_slv(opcode_type, 16#07#),
      1008 => to_slv(opcode_type, 16#09#),
      1009 => to_slv(opcode_type, 16#0B#),
      1010 => to_slv(opcode_type, 16#0D#),
      1011 => to_slv(opcode_type, 16#08#),
      1012 => to_slv(opcode_type, 16#0F#),
      1013 => to_slv(opcode_type, 16#0B#),
      1014 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#09#),
      1025 => to_slv(opcode_type, 16#02#),
      1026 => to_slv(opcode_type, 16#07#),
      1027 => to_slv(opcode_type, 16#01#),
      1028 => to_slv(opcode_type, 16#10#),
      1029 => to_slv(opcode_type, 16#03#),
      1030 => to_slv(opcode_type, 16#0F#),
      1031 => to_slv(opcode_type, 16#06#),
      1032 => to_slv(opcode_type, 16#08#),
      1033 => to_slv(opcode_type, 16#06#),
      1034 => to_slv(opcode_type, 16#11#),
      1035 => to_slv(opcode_type, 16#0B#),
      1036 => to_slv(opcode_type, 16#07#),
      1037 => to_slv(opcode_type, 16#0E#),
      1038 => to_slv(opcode_type, 16#0F#),
      1039 => to_slv(opcode_type, 16#07#),
      1040 => to_slv(opcode_type, 16#09#),
      1041 => to_slv(opcode_type, 16#CE#),
      1042 => to_slv(opcode_type, 16#0E#),
      1043 => to_slv(opcode_type, 16#06#),
      1044 => to_slv(opcode_type, 16#11#),
      1045 => to_slv(opcode_type, 16#0B#),
      1046 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#07#),
      1057 => to_slv(opcode_type, 16#09#),
      1058 => to_slv(opcode_type, 16#01#),
      1059 => to_slv(opcode_type, 16#03#),
      1060 => to_slv(opcode_type, 16#10#),
      1061 => to_slv(opcode_type, 16#06#),
      1062 => to_slv(opcode_type, 16#09#),
      1063 => to_slv(opcode_type, 16#11#),
      1064 => to_slv(opcode_type, 16#10#),
      1065 => to_slv(opcode_type, 16#05#),
      1066 => to_slv(opcode_type, 16#0E#),
      1067 => to_slv(opcode_type, 16#08#),
      1068 => to_slv(opcode_type, 16#06#),
      1069 => to_slv(opcode_type, 16#06#),
      1070 => to_slv(opcode_type, 16#11#),
      1071 => to_slv(opcode_type, 16#5A#),
      1072 => to_slv(opcode_type, 16#01#),
      1073 => to_slv(opcode_type, 16#0D#),
      1074 => to_slv(opcode_type, 16#02#),
      1075 => to_slv(opcode_type, 16#07#),
      1076 => to_slv(opcode_type, 16#0D#),
      1077 => to_slv(opcode_type, 16#0E#),
      1078 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#08#),
      1089 => to_slv(opcode_type, 16#08#),
      1090 => to_slv(opcode_type, 16#02#),
      1091 => to_slv(opcode_type, 16#05#),
      1092 => to_slv(opcode_type, 16#0F#),
      1093 => to_slv(opcode_type, 16#07#),
      1094 => to_slv(opcode_type, 16#02#),
      1095 => to_slv(opcode_type, 16#0D#),
      1096 => to_slv(opcode_type, 16#08#),
      1097 => to_slv(opcode_type, 16#0D#),
      1098 => to_slv(opcode_type, 16#0A#),
      1099 => to_slv(opcode_type, 16#09#),
      1100 => to_slv(opcode_type, 16#05#),
      1101 => to_slv(opcode_type, 16#09#),
      1102 => to_slv(opcode_type, 16#11#),
      1103 => to_slv(opcode_type, 16#0D#),
      1104 => to_slv(opcode_type, 16#06#),
      1105 => to_slv(opcode_type, 16#05#),
      1106 => to_slv(opcode_type, 16#0E#),
      1107 => to_slv(opcode_type, 16#07#),
      1108 => to_slv(opcode_type, 16#0F#),
      1109 => to_slv(opcode_type, 16#0F#),
      1110 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#08#),
      1121 => to_slv(opcode_type, 16#03#),
      1122 => to_slv(opcode_type, 16#07#),
      1123 => to_slv(opcode_type, 16#02#),
      1124 => to_slv(opcode_type, 16#0D#),
      1125 => to_slv(opcode_type, 16#05#),
      1126 => to_slv(opcode_type, 16#11#),
      1127 => to_slv(opcode_type, 16#09#),
      1128 => to_slv(opcode_type, 16#06#),
      1129 => to_slv(opcode_type, 16#06#),
      1130 => to_slv(opcode_type, 16#0D#),
      1131 => to_slv(opcode_type, 16#11#),
      1132 => to_slv(opcode_type, 16#07#),
      1133 => to_slv(opcode_type, 16#0E#),
      1134 => to_slv(opcode_type, 16#0D#),
      1135 => to_slv(opcode_type, 16#09#),
      1136 => to_slv(opcode_type, 16#07#),
      1137 => to_slv(opcode_type, 16#0B#),
      1138 => to_slv(opcode_type, 16#D4#),
      1139 => to_slv(opcode_type, 16#06#),
      1140 => to_slv(opcode_type, 16#11#),
      1141 => to_slv(opcode_type, 16#22#),
      1142 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#08#),
      1153 => to_slv(opcode_type, 16#04#),
      1154 => to_slv(opcode_type, 16#07#),
      1155 => to_slv(opcode_type, 16#03#),
      1156 => to_slv(opcode_type, 16#0F#),
      1157 => to_slv(opcode_type, 16#08#),
      1158 => to_slv(opcode_type, 16#E1#),
      1159 => to_slv(opcode_type, 16#0F#),
      1160 => to_slv(opcode_type, 16#08#),
      1161 => to_slv(opcode_type, 16#06#),
      1162 => to_slv(opcode_type, 16#08#),
      1163 => to_slv(opcode_type, 16#0D#),
      1164 => to_slv(opcode_type, 16#0D#),
      1165 => to_slv(opcode_type, 16#03#),
      1166 => to_slv(opcode_type, 16#11#),
      1167 => to_slv(opcode_type, 16#06#),
      1168 => to_slv(opcode_type, 16#08#),
      1169 => to_slv(opcode_type, 16#0B#),
      1170 => to_slv(opcode_type, 16#0A#),
      1171 => to_slv(opcode_type, 16#06#),
      1172 => to_slv(opcode_type, 16#B5#),
      1173 => to_slv(opcode_type, 16#11#),
      1174 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#06#),
      1185 => to_slv(opcode_type, 16#01#),
      1186 => to_slv(opcode_type, 16#09#),
      1187 => to_slv(opcode_type, 16#04#),
      1188 => to_slv(opcode_type, 16#11#),
      1189 => to_slv(opcode_type, 16#09#),
      1190 => to_slv(opcode_type, 16#0E#),
      1191 => to_slv(opcode_type, 16#10#),
      1192 => to_slv(opcode_type, 16#09#),
      1193 => to_slv(opcode_type, 16#07#),
      1194 => to_slv(opcode_type, 16#06#),
      1195 => to_slv(opcode_type, 16#8E#),
      1196 => to_slv(opcode_type, 16#0C#),
      1197 => to_slv(opcode_type, 16#06#),
      1198 => to_slv(opcode_type, 16#0A#),
      1199 => to_slv(opcode_type, 16#0D#),
      1200 => to_slv(opcode_type, 16#08#),
      1201 => to_slv(opcode_type, 16#03#),
      1202 => to_slv(opcode_type, 16#0D#),
      1203 => to_slv(opcode_type, 16#06#),
      1204 => to_slv(opcode_type, 16#10#),
      1205 => to_slv(opcode_type, 16#0C#),
      1206 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#06#),
      1217 => to_slv(opcode_type, 16#01#),
      1218 => to_slv(opcode_type, 16#09#),
      1219 => to_slv(opcode_type, 16#09#),
      1220 => to_slv(opcode_type, 16#11#),
      1221 => to_slv(opcode_type, 16#11#),
      1222 => to_slv(opcode_type, 16#09#),
      1223 => to_slv(opcode_type, 16#D8#),
      1224 => to_slv(opcode_type, 16#0C#),
      1225 => to_slv(opcode_type, 16#07#),
      1226 => to_slv(opcode_type, 16#08#),
      1227 => to_slv(opcode_type, 16#08#),
      1228 => to_slv(opcode_type, 16#0B#),
      1229 => to_slv(opcode_type, 16#0A#),
      1230 => to_slv(opcode_type, 16#02#),
      1231 => to_slv(opcode_type, 16#0C#),
      1232 => to_slv(opcode_type, 16#08#),
      1233 => to_slv(opcode_type, 16#02#),
      1234 => to_slv(opcode_type, 16#0E#),
      1235 => to_slv(opcode_type, 16#07#),
      1236 => to_slv(opcode_type, 16#0F#),
      1237 => to_slv(opcode_type, 16#0F#),
      1238 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#08#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#05#),
      1251 => to_slv(opcode_type, 16#04#),
      1252 => to_slv(opcode_type, 16#11#),
      1253 => to_slv(opcode_type, 16#04#),
      1254 => to_slv(opcode_type, 16#04#),
      1255 => to_slv(opcode_type, 16#0D#),
      1256 => to_slv(opcode_type, 16#09#),
      1257 => to_slv(opcode_type, 16#06#),
      1258 => to_slv(opcode_type, 16#07#),
      1259 => to_slv(opcode_type, 16#0A#),
      1260 => to_slv(opcode_type, 16#10#),
      1261 => to_slv(opcode_type, 16#05#),
      1262 => to_slv(opcode_type, 16#0C#),
      1263 => to_slv(opcode_type, 16#07#),
      1264 => to_slv(opcode_type, 16#06#),
      1265 => to_slv(opcode_type, 16#0C#),
      1266 => to_slv(opcode_type, 16#0C#),
      1267 => to_slv(opcode_type, 16#08#),
      1268 => to_slv(opcode_type, 16#D1#),
      1269 => to_slv(opcode_type, 16#11#),
      1270 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#08#),
      1281 => to_slv(opcode_type, 16#02#),
      1282 => to_slv(opcode_type, 16#06#),
      1283 => to_slv(opcode_type, 16#03#),
      1284 => to_slv(opcode_type, 16#0B#),
      1285 => to_slv(opcode_type, 16#08#),
      1286 => to_slv(opcode_type, 16#11#),
      1287 => to_slv(opcode_type, 16#0B#),
      1288 => to_slv(opcode_type, 16#09#),
      1289 => to_slv(opcode_type, 16#09#),
      1290 => to_slv(opcode_type, 16#01#),
      1291 => to_slv(opcode_type, 16#13#),
      1292 => to_slv(opcode_type, 16#06#),
      1293 => to_slv(opcode_type, 16#0C#),
      1294 => to_slv(opcode_type, 16#0F#),
      1295 => to_slv(opcode_type, 16#06#),
      1296 => to_slv(opcode_type, 16#09#),
      1297 => to_slv(opcode_type, 16#0A#),
      1298 => to_slv(opcode_type, 16#0D#),
      1299 => to_slv(opcode_type, 16#07#),
      1300 => to_slv(opcode_type, 16#0D#),
      1301 => to_slv(opcode_type, 16#0B#),
      1302 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#07#),
      1313 => to_slv(opcode_type, 16#04#),
      1314 => to_slv(opcode_type, 16#08#),
      1315 => to_slv(opcode_type, 16#03#),
      1316 => to_slv(opcode_type, 16#0C#),
      1317 => to_slv(opcode_type, 16#05#),
      1318 => to_slv(opcode_type, 16#0E#),
      1319 => to_slv(opcode_type, 16#09#),
      1320 => to_slv(opcode_type, 16#08#),
      1321 => to_slv(opcode_type, 16#06#),
      1322 => to_slv(opcode_type, 16#10#),
      1323 => to_slv(opcode_type, 16#11#),
      1324 => to_slv(opcode_type, 16#06#),
      1325 => to_slv(opcode_type, 16#0B#),
      1326 => to_slv(opcode_type, 16#0F#),
      1327 => to_slv(opcode_type, 16#07#),
      1328 => to_slv(opcode_type, 16#07#),
      1329 => to_slv(opcode_type, 16#27#),
      1330 => to_slv(opcode_type, 16#11#),
      1331 => to_slv(opcode_type, 16#09#),
      1332 => to_slv(opcode_type, 16#0B#),
      1333 => to_slv(opcode_type, 16#0A#),
      1334 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#07#),
      1345 => to_slv(opcode_type, 16#07#),
      1346 => to_slv(opcode_type, 16#01#),
      1347 => to_slv(opcode_type, 16#03#),
      1348 => to_slv(opcode_type, 16#0A#),
      1349 => to_slv(opcode_type, 16#02#),
      1350 => to_slv(opcode_type, 16#02#),
      1351 => to_slv(opcode_type, 16#0A#),
      1352 => to_slv(opcode_type, 16#09#),
      1353 => to_slv(opcode_type, 16#07#),
      1354 => to_slv(opcode_type, 16#08#),
      1355 => to_slv(opcode_type, 16#B1#),
      1356 => to_slv(opcode_type, 16#0F#),
      1357 => to_slv(opcode_type, 16#04#),
      1358 => to_slv(opcode_type, 16#0D#),
      1359 => to_slv(opcode_type, 16#06#),
      1360 => to_slv(opcode_type, 16#08#),
      1361 => to_slv(opcode_type, 16#0C#),
      1362 => to_slv(opcode_type, 16#11#),
      1363 => to_slv(opcode_type, 16#09#),
      1364 => to_slv(opcode_type, 16#10#),
      1365 => to_slv(opcode_type, 16#0B#),
      1366 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#09#),
      1377 => to_slv(opcode_type, 16#02#),
      1378 => to_slv(opcode_type, 16#06#),
      1379 => to_slv(opcode_type, 16#03#),
      1380 => to_slv(opcode_type, 16#DF#),
      1381 => to_slv(opcode_type, 16#05#),
      1382 => to_slv(opcode_type, 16#BE#),
      1383 => to_slv(opcode_type, 16#06#),
      1384 => to_slv(opcode_type, 16#08#),
      1385 => to_slv(opcode_type, 16#09#),
      1386 => to_slv(opcode_type, 16#0F#),
      1387 => to_slv(opcode_type, 16#0E#),
      1388 => to_slv(opcode_type, 16#08#),
      1389 => to_slv(opcode_type, 16#20#),
      1390 => to_slv(opcode_type, 16#0D#),
      1391 => to_slv(opcode_type, 16#06#),
      1392 => to_slv(opcode_type, 16#07#),
      1393 => to_slv(opcode_type, 16#0F#),
      1394 => to_slv(opcode_type, 16#10#),
      1395 => to_slv(opcode_type, 16#06#),
      1396 => to_slv(opcode_type, 16#0C#),
      1397 => to_slv(opcode_type, 16#0A#),
      1398 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#05#),
      1410 => to_slv(opcode_type, 16#09#),
      1411 => to_slv(opcode_type, 16#04#),
      1412 => to_slv(opcode_type, 16#0B#),
      1413 => to_slv(opcode_type, 16#08#),
      1414 => to_slv(opcode_type, 16#0F#),
      1415 => to_slv(opcode_type, 16#11#),
      1416 => to_slv(opcode_type, 16#09#),
      1417 => to_slv(opcode_type, 16#09#),
      1418 => to_slv(opcode_type, 16#09#),
      1419 => to_slv(opcode_type, 16#0D#),
      1420 => to_slv(opcode_type, 16#0F#),
      1421 => to_slv(opcode_type, 16#09#),
      1422 => to_slv(opcode_type, 16#0E#),
      1423 => to_slv(opcode_type, 16#54#),
      1424 => to_slv(opcode_type, 16#06#),
      1425 => to_slv(opcode_type, 16#07#),
      1426 => to_slv(opcode_type, 16#0A#),
      1427 => to_slv(opcode_type, 16#0C#),
      1428 => to_slv(opcode_type, 16#03#),
      1429 => to_slv(opcode_type, 16#A0#),
      1430 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#09#),
      1441 => to_slv(opcode_type, 16#07#),
      1442 => to_slv(opcode_type, 16#03#),
      1443 => to_slv(opcode_type, 16#02#),
      1444 => to_slv(opcode_type, 16#0F#),
      1445 => to_slv(opcode_type, 16#03#),
      1446 => to_slv(opcode_type, 16#08#),
      1447 => to_slv(opcode_type, 16#0F#),
      1448 => to_slv(opcode_type, 16#0A#),
      1449 => to_slv(opcode_type, 16#06#),
      1450 => to_slv(opcode_type, 16#06#),
      1451 => to_slv(opcode_type, 16#07#),
      1452 => to_slv(opcode_type, 16#0F#),
      1453 => to_slv(opcode_type, 16#10#),
      1454 => to_slv(opcode_type, 16#05#),
      1455 => to_slv(opcode_type, 16#11#),
      1456 => to_slv(opcode_type, 16#09#),
      1457 => to_slv(opcode_type, 16#01#),
      1458 => to_slv(opcode_type, 16#0C#),
      1459 => to_slv(opcode_type, 16#07#),
      1460 => to_slv(opcode_type, 16#0B#),
      1461 => to_slv(opcode_type, 16#0D#),
      1462 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#08#),
      1473 => to_slv(opcode_type, 16#07#),
      1474 => to_slv(opcode_type, 16#08#),
      1475 => to_slv(opcode_type, 16#09#),
      1476 => to_slv(opcode_type, 16#0E#),
      1477 => to_slv(opcode_type, 16#0D#),
      1478 => to_slv(opcode_type, 16#01#),
      1479 => to_slv(opcode_type, 16#0F#),
      1480 => to_slv(opcode_type, 16#07#),
      1481 => to_slv(opcode_type, 16#04#),
      1482 => to_slv(opcode_type, 16#0D#),
      1483 => to_slv(opcode_type, 16#02#),
      1484 => to_slv(opcode_type, 16#0A#),
      1485 => to_slv(opcode_type, 16#09#),
      1486 => to_slv(opcode_type, 16#01#),
      1487 => to_slv(opcode_type, 16#08#),
      1488 => to_slv(opcode_type, 16#11#),
      1489 => to_slv(opcode_type, 16#0E#),
      1490 => to_slv(opcode_type, 16#09#),
      1491 => to_slv(opcode_type, 16#03#),
      1492 => to_slv(opcode_type, 16#0A#),
      1493 => to_slv(opcode_type, 16#0A#),
      1494 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#09#),
      1505 => to_slv(opcode_type, 16#04#),
      1506 => to_slv(opcode_type, 16#07#),
      1507 => to_slv(opcode_type, 16#07#),
      1508 => to_slv(opcode_type, 16#7D#),
      1509 => to_slv(opcode_type, 16#0B#),
      1510 => to_slv(opcode_type, 16#07#),
      1511 => to_slv(opcode_type, 16#0F#),
      1512 => to_slv(opcode_type, 16#10#),
      1513 => to_slv(opcode_type, 16#07#),
      1514 => to_slv(opcode_type, 16#08#),
      1515 => to_slv(opcode_type, 16#05#),
      1516 => to_slv(opcode_type, 16#0C#),
      1517 => to_slv(opcode_type, 16#01#),
      1518 => to_slv(opcode_type, 16#0C#),
      1519 => to_slv(opcode_type, 16#09#),
      1520 => to_slv(opcode_type, 16#08#),
      1521 => to_slv(opcode_type, 16#11#),
      1522 => to_slv(opcode_type, 16#11#),
      1523 => to_slv(opcode_type, 16#06#),
      1524 => to_slv(opcode_type, 16#11#),
      1525 => to_slv(opcode_type, 16#0C#),
      1526 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#08#),
      1537 => to_slv(opcode_type, 16#04#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#06#),
      1540 => to_slv(opcode_type, 16#11#),
      1541 => to_slv(opcode_type, 16#0C#),
      1542 => to_slv(opcode_type, 16#05#),
      1543 => to_slv(opcode_type, 16#0C#),
      1544 => to_slv(opcode_type, 16#09#),
      1545 => to_slv(opcode_type, 16#08#),
      1546 => to_slv(opcode_type, 16#07#),
      1547 => to_slv(opcode_type, 16#0B#),
      1548 => to_slv(opcode_type, 16#0A#),
      1549 => to_slv(opcode_type, 16#07#),
      1550 => to_slv(opcode_type, 16#0A#),
      1551 => to_slv(opcode_type, 16#0D#),
      1552 => to_slv(opcode_type, 16#08#),
      1553 => to_slv(opcode_type, 16#09#),
      1554 => to_slv(opcode_type, 16#0F#),
      1555 => to_slv(opcode_type, 16#33#),
      1556 => to_slv(opcode_type, 16#01#),
      1557 => to_slv(opcode_type, 16#11#),
      1558 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#06#),
      1569 => to_slv(opcode_type, 16#05#),
      1570 => to_slv(opcode_type, 16#07#),
      1571 => to_slv(opcode_type, 16#09#),
      1572 => to_slv(opcode_type, 16#10#),
      1573 => to_slv(opcode_type, 16#0C#),
      1574 => to_slv(opcode_type, 16#04#),
      1575 => to_slv(opcode_type, 16#0F#),
      1576 => to_slv(opcode_type, 16#09#),
      1577 => to_slv(opcode_type, 16#06#),
      1578 => to_slv(opcode_type, 16#02#),
      1579 => to_slv(opcode_type, 16#0C#),
      1580 => to_slv(opcode_type, 16#06#),
      1581 => to_slv(opcode_type, 16#0A#),
      1582 => to_slv(opcode_type, 16#0A#),
      1583 => to_slv(opcode_type, 16#06#),
      1584 => to_slv(opcode_type, 16#06#),
      1585 => to_slv(opcode_type, 16#10#),
      1586 => to_slv(opcode_type, 16#0F#),
      1587 => to_slv(opcode_type, 16#06#),
      1588 => to_slv(opcode_type, 16#11#),
      1589 => to_slv(opcode_type, 16#0D#),
      1590 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#02#),
      1602 => to_slv(opcode_type, 16#07#),
      1603 => to_slv(opcode_type, 16#03#),
      1604 => to_slv(opcode_type, 16#0B#),
      1605 => to_slv(opcode_type, 16#03#),
      1606 => to_slv(opcode_type, 16#0D#),
      1607 => to_slv(opcode_type, 16#07#),
      1608 => to_slv(opcode_type, 16#09#),
      1609 => to_slv(opcode_type, 16#08#),
      1610 => to_slv(opcode_type, 16#0C#),
      1611 => to_slv(opcode_type, 16#0A#),
      1612 => to_slv(opcode_type, 16#09#),
      1613 => to_slv(opcode_type, 16#0F#),
      1614 => to_slv(opcode_type, 16#0E#),
      1615 => to_slv(opcode_type, 16#06#),
      1616 => to_slv(opcode_type, 16#06#),
      1617 => to_slv(opcode_type, 16#0B#),
      1618 => to_slv(opcode_type, 16#10#),
      1619 => to_slv(opcode_type, 16#09#),
      1620 => to_slv(opcode_type, 16#11#),
      1621 => to_slv(opcode_type, 16#0B#),
      1622 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#09#),
      1633 => to_slv(opcode_type, 16#09#),
      1634 => to_slv(opcode_type, 16#07#),
      1635 => to_slv(opcode_type, 16#06#),
      1636 => to_slv(opcode_type, 16#0A#),
      1637 => to_slv(opcode_type, 16#10#),
      1638 => to_slv(opcode_type, 16#07#),
      1639 => to_slv(opcode_type, 16#0C#),
      1640 => to_slv(opcode_type, 16#0A#),
      1641 => to_slv(opcode_type, 16#07#),
      1642 => to_slv(opcode_type, 16#05#),
      1643 => to_slv(opcode_type, 16#59#),
      1644 => to_slv(opcode_type, 16#02#),
      1645 => to_slv(opcode_type, 16#0B#),
      1646 => to_slv(opcode_type, 16#03#),
      1647 => to_slv(opcode_type, 16#07#),
      1648 => to_slv(opcode_type, 16#08#),
      1649 => to_slv(opcode_type, 16#0B#),
      1650 => to_slv(opcode_type, 16#11#),
      1651 => to_slv(opcode_type, 16#07#),
      1652 => to_slv(opcode_type, 16#10#),
      1653 => to_slv(opcode_type, 16#0C#),
      1654 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#06#),
      1665 => to_slv(opcode_type, 16#03#),
      1666 => to_slv(opcode_type, 16#08#),
      1667 => to_slv(opcode_type, 16#07#),
      1668 => to_slv(opcode_type, 16#8B#),
      1669 => to_slv(opcode_type, 16#39#),
      1670 => to_slv(opcode_type, 16#01#),
      1671 => to_slv(opcode_type, 16#11#),
      1672 => to_slv(opcode_type, 16#07#),
      1673 => to_slv(opcode_type, 16#08#),
      1674 => to_slv(opcode_type, 16#07#),
      1675 => to_slv(opcode_type, 16#0E#),
      1676 => to_slv(opcode_type, 16#10#),
      1677 => to_slv(opcode_type, 16#03#),
      1678 => to_slv(opcode_type, 16#0C#),
      1679 => to_slv(opcode_type, 16#08#),
      1680 => to_slv(opcode_type, 16#09#),
      1681 => to_slv(opcode_type, 16#0C#),
      1682 => to_slv(opcode_type, 16#0A#),
      1683 => to_slv(opcode_type, 16#08#),
      1684 => to_slv(opcode_type, 16#0B#),
      1685 => to_slv(opcode_type, 16#11#),
      1686 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#09#),
      1697 => to_slv(opcode_type, 16#04#),
      1698 => to_slv(opcode_type, 16#07#),
      1699 => to_slv(opcode_type, 16#07#),
      1700 => to_slv(opcode_type, 16#10#),
      1701 => to_slv(opcode_type, 16#D4#),
      1702 => to_slv(opcode_type, 16#07#),
      1703 => to_slv(opcode_type, 16#0E#),
      1704 => to_slv(opcode_type, 16#0B#),
      1705 => to_slv(opcode_type, 16#09#),
      1706 => to_slv(opcode_type, 16#09#),
      1707 => to_slv(opcode_type, 16#07#),
      1708 => to_slv(opcode_type, 16#0F#),
      1709 => to_slv(opcode_type, 16#0E#),
      1710 => to_slv(opcode_type, 16#06#),
      1711 => to_slv(opcode_type, 16#0A#),
      1712 => to_slv(opcode_type, 16#0D#),
      1713 => to_slv(opcode_type, 16#09#),
      1714 => to_slv(opcode_type, 16#06#),
      1715 => to_slv(opcode_type, 16#0C#),
      1716 => to_slv(opcode_type, 16#0C#),
      1717 => to_slv(opcode_type, 16#10#),
      1718 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#07#),
      1729 => to_slv(opcode_type, 16#09#),
      1730 => to_slv(opcode_type, 16#01#),
      1731 => to_slv(opcode_type, 16#01#),
      1732 => to_slv(opcode_type, 16#0E#),
      1733 => to_slv(opcode_type, 16#05#),
      1734 => to_slv(opcode_type, 16#09#),
      1735 => to_slv(opcode_type, 16#0B#),
      1736 => to_slv(opcode_type, 16#0C#),
      1737 => to_slv(opcode_type, 16#06#),
      1738 => to_slv(opcode_type, 16#09#),
      1739 => to_slv(opcode_type, 16#06#),
      1740 => to_slv(opcode_type, 16#0B#),
      1741 => to_slv(opcode_type, 16#0E#),
      1742 => to_slv(opcode_type, 16#06#),
      1743 => to_slv(opcode_type, 16#0E#),
      1744 => to_slv(opcode_type, 16#0C#),
      1745 => to_slv(opcode_type, 16#08#),
      1746 => to_slv(opcode_type, 16#07#),
      1747 => to_slv(opcode_type, 16#10#),
      1748 => to_slv(opcode_type, 16#0E#),
      1749 => to_slv(opcode_type, 16#0B#),
      1750 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#08#),
      1761 => to_slv(opcode_type, 16#02#),
      1762 => to_slv(opcode_type, 16#06#),
      1763 => to_slv(opcode_type, 16#04#),
      1764 => to_slv(opcode_type, 16#0B#),
      1765 => to_slv(opcode_type, 16#01#),
      1766 => to_slv(opcode_type, 16#0A#),
      1767 => to_slv(opcode_type, 16#07#),
      1768 => to_slv(opcode_type, 16#09#),
      1769 => to_slv(opcode_type, 16#09#),
      1770 => to_slv(opcode_type, 16#0C#),
      1771 => to_slv(opcode_type, 16#0D#),
      1772 => to_slv(opcode_type, 16#07#),
      1773 => to_slv(opcode_type, 16#0D#),
      1774 => to_slv(opcode_type, 16#0C#),
      1775 => to_slv(opcode_type, 16#09#),
      1776 => to_slv(opcode_type, 16#08#),
      1777 => to_slv(opcode_type, 16#0E#),
      1778 => to_slv(opcode_type, 16#0A#),
      1779 => to_slv(opcode_type, 16#06#),
      1780 => to_slv(opcode_type, 16#0C#),
      1781 => to_slv(opcode_type, 16#11#),
      1782 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#08#),
      1793 => to_slv(opcode_type, 16#07#),
      1794 => to_slv(opcode_type, 16#03#),
      1795 => to_slv(opcode_type, 16#09#),
      1796 => to_slv(opcode_type, 16#0B#),
      1797 => to_slv(opcode_type, 16#11#),
      1798 => to_slv(opcode_type, 16#06#),
      1799 => to_slv(opcode_type, 16#08#),
      1800 => to_slv(opcode_type, 16#11#),
      1801 => to_slv(opcode_type, 16#0B#),
      1802 => to_slv(opcode_type, 16#05#),
      1803 => to_slv(opcode_type, 16#0C#),
      1804 => to_slv(opcode_type, 16#08#),
      1805 => to_slv(opcode_type, 16#06#),
      1806 => to_slv(opcode_type, 16#03#),
      1807 => to_slv(opcode_type, 16#B8#),
      1808 => to_slv(opcode_type, 16#06#),
      1809 => to_slv(opcode_type, 16#0B#),
      1810 => to_slv(opcode_type, 16#0B#),
      1811 => to_slv(opcode_type, 16#04#),
      1812 => to_slv(opcode_type, 16#05#),
      1813 => to_slv(opcode_type, 16#0A#),
      1814 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#07#),
      1825 => to_slv(opcode_type, 16#07#),
      1826 => to_slv(opcode_type, 16#02#),
      1827 => to_slv(opcode_type, 16#04#),
      1828 => to_slv(opcode_type, 16#0C#),
      1829 => to_slv(opcode_type, 16#03#),
      1830 => to_slv(opcode_type, 16#04#),
      1831 => to_slv(opcode_type, 16#0E#),
      1832 => to_slv(opcode_type, 16#07#),
      1833 => to_slv(opcode_type, 16#09#),
      1834 => to_slv(opcode_type, 16#04#),
      1835 => to_slv(opcode_type, 16#0E#),
      1836 => to_slv(opcode_type, 16#08#),
      1837 => to_slv(opcode_type, 16#0C#),
      1838 => to_slv(opcode_type, 16#0C#),
      1839 => to_slv(opcode_type, 16#07#),
      1840 => to_slv(opcode_type, 16#06#),
      1841 => to_slv(opcode_type, 16#0C#),
      1842 => to_slv(opcode_type, 16#0A#),
      1843 => to_slv(opcode_type, 16#08#),
      1844 => to_slv(opcode_type, 16#0D#),
      1845 => to_slv(opcode_type, 16#0E#),
      1846 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#09#),
      1857 => to_slv(opcode_type, 16#04#),
      1858 => to_slv(opcode_type, 16#07#),
      1859 => to_slv(opcode_type, 16#02#),
      1860 => to_slv(opcode_type, 16#0D#),
      1861 => to_slv(opcode_type, 16#07#),
      1862 => to_slv(opcode_type, 16#5A#),
      1863 => to_slv(opcode_type, 16#11#),
      1864 => to_slv(opcode_type, 16#06#),
      1865 => to_slv(opcode_type, 16#09#),
      1866 => to_slv(opcode_type, 16#05#),
      1867 => to_slv(opcode_type, 16#AD#),
      1868 => to_slv(opcode_type, 16#06#),
      1869 => to_slv(opcode_type, 16#0B#),
      1870 => to_slv(opcode_type, 16#0D#),
      1871 => to_slv(opcode_type, 16#09#),
      1872 => to_slv(opcode_type, 16#07#),
      1873 => to_slv(opcode_type, 16#8F#),
      1874 => to_slv(opcode_type, 16#0B#),
      1875 => to_slv(opcode_type, 16#08#),
      1876 => to_slv(opcode_type, 16#10#),
      1877 => to_slv(opcode_type, 16#0F#),
      1878 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#08#),
      1889 => to_slv(opcode_type, 16#07#),
      1890 => to_slv(opcode_type, 16#06#),
      1891 => to_slv(opcode_type, 16#02#),
      1892 => to_slv(opcode_type, 16#0D#),
      1893 => to_slv(opcode_type, 16#05#),
      1894 => to_slv(opcode_type, 16#0B#),
      1895 => to_slv(opcode_type, 16#05#),
      1896 => to_slv(opcode_type, 16#09#),
      1897 => to_slv(opcode_type, 16#7B#),
      1898 => to_slv(opcode_type, 16#10#),
      1899 => to_slv(opcode_type, 16#09#),
      1900 => to_slv(opcode_type, 16#04#),
      1901 => to_slv(opcode_type, 16#08#),
      1902 => to_slv(opcode_type, 16#0A#),
      1903 => to_slv(opcode_type, 16#FF#),
      1904 => to_slv(opcode_type, 16#08#),
      1905 => to_slv(opcode_type, 16#08#),
      1906 => to_slv(opcode_type, 16#11#),
      1907 => to_slv(opcode_type, 16#0A#),
      1908 => to_slv(opcode_type, 16#03#),
      1909 => to_slv(opcode_type, 16#0D#),
      1910 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#08#),
      1921 => to_slv(opcode_type, 16#03#),
      1922 => to_slv(opcode_type, 16#06#),
      1923 => to_slv(opcode_type, 16#06#),
      1924 => to_slv(opcode_type, 16#D2#),
      1925 => to_slv(opcode_type, 16#E1#),
      1926 => to_slv(opcode_type, 16#04#),
      1927 => to_slv(opcode_type, 16#11#),
      1928 => to_slv(opcode_type, 16#09#),
      1929 => to_slv(opcode_type, 16#08#),
      1930 => to_slv(opcode_type, 16#04#),
      1931 => to_slv(opcode_type, 16#0C#),
      1932 => to_slv(opcode_type, 16#08#),
      1933 => to_slv(opcode_type, 16#10#),
      1934 => to_slv(opcode_type, 16#0A#),
      1935 => to_slv(opcode_type, 16#09#),
      1936 => to_slv(opcode_type, 16#06#),
      1937 => to_slv(opcode_type, 16#0D#),
      1938 => to_slv(opcode_type, 16#0A#),
      1939 => to_slv(opcode_type, 16#09#),
      1940 => to_slv(opcode_type, 16#C1#),
      1941 => to_slv(opcode_type, 16#0A#),
      1942 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#07#),
      1953 => to_slv(opcode_type, 16#07#),
      1954 => to_slv(opcode_type, 16#07#),
      1955 => to_slv(opcode_type, 16#02#),
      1956 => to_slv(opcode_type, 16#0E#),
      1957 => to_slv(opcode_type, 16#08#),
      1958 => to_slv(opcode_type, 16#0A#),
      1959 => to_slv(opcode_type, 16#77#),
      1960 => to_slv(opcode_type, 16#02#),
      1961 => to_slv(opcode_type, 16#08#),
      1962 => to_slv(opcode_type, 16#0D#),
      1963 => to_slv(opcode_type, 16#19#),
      1964 => to_slv(opcode_type, 16#08#),
      1965 => to_slv(opcode_type, 16#04#),
      1966 => to_slv(opcode_type, 16#04#),
      1967 => to_slv(opcode_type, 16#11#),
      1968 => to_slv(opcode_type, 16#08#),
      1969 => to_slv(opcode_type, 16#06#),
      1970 => to_slv(opcode_type, 16#0E#),
      1971 => to_slv(opcode_type, 16#0F#),
      1972 => to_slv(opcode_type, 16#02#),
      1973 => to_slv(opcode_type, 16#10#),
      1974 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#08#),
      1985 => to_slv(opcode_type, 16#07#),
      1986 => to_slv(opcode_type, 16#08#),
      1987 => to_slv(opcode_type, 16#05#),
      1988 => to_slv(opcode_type, 16#0C#),
      1989 => to_slv(opcode_type, 16#03#),
      1990 => to_slv(opcode_type, 16#0F#),
      1991 => to_slv(opcode_type, 16#05#),
      1992 => to_slv(opcode_type, 16#05#),
      1993 => to_slv(opcode_type, 16#11#),
      1994 => to_slv(opcode_type, 16#09#),
      1995 => to_slv(opcode_type, 16#08#),
      1996 => to_slv(opcode_type, 16#05#),
      1997 => to_slv(opcode_type, 16#11#),
      1998 => to_slv(opcode_type, 16#05#),
      1999 => to_slv(opcode_type, 16#10#),
      2000 => to_slv(opcode_type, 16#06#),
      2001 => to_slv(opcode_type, 16#06#),
      2002 => to_slv(opcode_type, 16#11#),
      2003 => to_slv(opcode_type, 16#0F#),
      2004 => to_slv(opcode_type, 16#04#),
      2005 => to_slv(opcode_type, 16#0B#),
      2006 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#08#),
      2017 => to_slv(opcode_type, 16#02#),
      2018 => to_slv(opcode_type, 16#08#),
      2019 => to_slv(opcode_type, 16#07#),
      2020 => to_slv(opcode_type, 16#0A#),
      2021 => to_slv(opcode_type, 16#0C#),
      2022 => to_slv(opcode_type, 16#08#),
      2023 => to_slv(opcode_type, 16#10#),
      2024 => to_slv(opcode_type, 16#0E#),
      2025 => to_slv(opcode_type, 16#07#),
      2026 => to_slv(opcode_type, 16#09#),
      2027 => to_slv(opcode_type, 16#06#),
      2028 => to_slv(opcode_type, 16#0F#),
      2029 => to_slv(opcode_type, 16#10#),
      2030 => to_slv(opcode_type, 16#07#),
      2031 => to_slv(opcode_type, 16#0D#),
      2032 => to_slv(opcode_type, 16#10#),
      2033 => to_slv(opcode_type, 16#09#),
      2034 => to_slv(opcode_type, 16#08#),
      2035 => to_slv(opcode_type, 16#0D#),
      2036 => to_slv(opcode_type, 16#0D#),
      2037 => to_slv(opcode_type, 16#0B#),
      2038 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#07#),
      2049 => to_slv(opcode_type, 16#02#),
      2050 => to_slv(opcode_type, 16#09#),
      2051 => to_slv(opcode_type, 16#05#),
      2052 => to_slv(opcode_type, 16#0C#),
      2053 => to_slv(opcode_type, 16#09#),
      2054 => to_slv(opcode_type, 16#11#),
      2055 => to_slv(opcode_type, 16#0F#),
      2056 => to_slv(opcode_type, 16#07#),
      2057 => to_slv(opcode_type, 16#08#),
      2058 => to_slv(opcode_type, 16#01#),
      2059 => to_slv(opcode_type, 16#10#),
      2060 => to_slv(opcode_type, 16#09#),
      2061 => to_slv(opcode_type, 16#0E#),
      2062 => to_slv(opcode_type, 16#0C#),
      2063 => to_slv(opcode_type, 16#09#),
      2064 => to_slv(opcode_type, 16#07#),
      2065 => to_slv(opcode_type, 16#0E#),
      2066 => to_slv(opcode_type, 16#0E#),
      2067 => to_slv(opcode_type, 16#08#),
      2068 => to_slv(opcode_type, 16#10#),
      2069 => to_slv(opcode_type, 16#0B#),
      2070 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#06#),
      2081 => to_slv(opcode_type, 16#02#),
      2082 => to_slv(opcode_type, 16#07#),
      2083 => to_slv(opcode_type, 16#09#),
      2084 => to_slv(opcode_type, 16#0F#),
      2085 => to_slv(opcode_type, 16#0E#),
      2086 => to_slv(opcode_type, 16#05#),
      2087 => to_slv(opcode_type, 16#0F#),
      2088 => to_slv(opcode_type, 16#08#),
      2089 => to_slv(opcode_type, 16#09#),
      2090 => to_slv(opcode_type, 16#01#),
      2091 => to_slv(opcode_type, 16#0A#),
      2092 => to_slv(opcode_type, 16#06#),
      2093 => to_slv(opcode_type, 16#11#),
      2094 => to_slv(opcode_type, 16#0E#),
      2095 => to_slv(opcode_type, 16#06#),
      2096 => to_slv(opcode_type, 16#07#),
      2097 => to_slv(opcode_type, 16#0F#),
      2098 => to_slv(opcode_type, 16#0D#),
      2099 => to_slv(opcode_type, 16#09#),
      2100 => to_slv(opcode_type, 16#0A#),
      2101 => to_slv(opcode_type, 16#0F#),
      2102 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#06#),
      2113 => to_slv(opcode_type, 16#07#),
      2114 => to_slv(opcode_type, 16#03#),
      2115 => to_slv(opcode_type, 16#05#),
      2116 => to_slv(opcode_type, 16#0A#),
      2117 => to_slv(opcode_type, 16#01#),
      2118 => to_slv(opcode_type, 16#04#),
      2119 => to_slv(opcode_type, 16#0C#),
      2120 => to_slv(opcode_type, 16#06#),
      2121 => to_slv(opcode_type, 16#09#),
      2122 => to_slv(opcode_type, 16#06#),
      2123 => to_slv(opcode_type, 16#10#),
      2124 => to_slv(opcode_type, 16#0E#),
      2125 => to_slv(opcode_type, 16#07#),
      2126 => to_slv(opcode_type, 16#0C#),
      2127 => to_slv(opcode_type, 16#0B#),
      2128 => to_slv(opcode_type, 16#09#),
      2129 => to_slv(opcode_type, 16#05#),
      2130 => to_slv(opcode_type, 16#11#),
      2131 => to_slv(opcode_type, 16#06#),
      2132 => to_slv(opcode_type, 16#0C#),
      2133 => to_slv(opcode_type, 16#0E#),
      2134 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#06#),
      2145 => to_slv(opcode_type, 16#02#),
      2146 => to_slv(opcode_type, 16#08#),
      2147 => to_slv(opcode_type, 16#02#),
      2148 => to_slv(opcode_type, 16#C4#),
      2149 => to_slv(opcode_type, 16#06#),
      2150 => to_slv(opcode_type, 16#0C#),
      2151 => to_slv(opcode_type, 16#0B#),
      2152 => to_slv(opcode_type, 16#09#),
      2153 => to_slv(opcode_type, 16#09#),
      2154 => to_slv(opcode_type, 16#07#),
      2155 => to_slv(opcode_type, 16#0B#),
      2156 => to_slv(opcode_type, 16#11#),
      2157 => to_slv(opcode_type, 16#01#),
      2158 => to_slv(opcode_type, 16#0A#),
      2159 => to_slv(opcode_type, 16#07#),
      2160 => to_slv(opcode_type, 16#08#),
      2161 => to_slv(opcode_type, 16#0C#),
      2162 => to_slv(opcode_type, 16#7B#),
      2163 => to_slv(opcode_type, 16#06#),
      2164 => to_slv(opcode_type, 16#10#),
      2165 => to_slv(opcode_type, 16#0B#),
      2166 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#07#),
      2177 => to_slv(opcode_type, 16#03#),
      2178 => to_slv(opcode_type, 16#09#),
      2179 => to_slv(opcode_type, 16#03#),
      2180 => to_slv(opcode_type, 16#0C#),
      2181 => to_slv(opcode_type, 16#03#),
      2182 => to_slv(opcode_type, 16#0C#),
      2183 => to_slv(opcode_type, 16#08#),
      2184 => to_slv(opcode_type, 16#09#),
      2185 => to_slv(opcode_type, 16#09#),
      2186 => to_slv(opcode_type, 16#0D#),
      2187 => to_slv(opcode_type, 16#0E#),
      2188 => to_slv(opcode_type, 16#09#),
      2189 => to_slv(opcode_type, 16#0D#),
      2190 => to_slv(opcode_type, 16#10#),
      2191 => to_slv(opcode_type, 16#06#),
      2192 => to_slv(opcode_type, 16#08#),
      2193 => to_slv(opcode_type, 16#0F#),
      2194 => to_slv(opcode_type, 16#11#),
      2195 => to_slv(opcode_type, 16#08#),
      2196 => to_slv(opcode_type, 16#0F#),
      2197 => to_slv(opcode_type, 16#10#),
      2198 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#09#),
      2209 => to_slv(opcode_type, 16#08#),
      2210 => to_slv(opcode_type, 16#07#),
      2211 => to_slv(opcode_type, 16#02#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#06#),
      2214 => to_slv(opcode_type, 16#0F#),
      2215 => to_slv(opcode_type, 16#10#),
      2216 => to_slv(opcode_type, 16#01#),
      2217 => to_slv(opcode_type, 16#03#),
      2218 => to_slv(opcode_type, 16#0B#),
      2219 => to_slv(opcode_type, 16#07#),
      2220 => to_slv(opcode_type, 16#02#),
      2221 => to_slv(opcode_type, 16#04#),
      2222 => to_slv(opcode_type, 16#11#),
      2223 => to_slv(opcode_type, 16#07#),
      2224 => to_slv(opcode_type, 16#06#),
      2225 => to_slv(opcode_type, 16#0C#),
      2226 => to_slv(opcode_type, 16#0A#),
      2227 => to_slv(opcode_type, 16#08#),
      2228 => to_slv(opcode_type, 16#0E#),
      2229 => to_slv(opcode_type, 16#0D#),
      2230 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#09#),
      2241 => to_slv(opcode_type, 16#04#),
      2242 => to_slv(opcode_type, 16#06#),
      2243 => to_slv(opcode_type, 16#03#),
      2244 => to_slv(opcode_type, 16#0E#),
      2245 => to_slv(opcode_type, 16#07#),
      2246 => to_slv(opcode_type, 16#0D#),
      2247 => to_slv(opcode_type, 16#0B#),
      2248 => to_slv(opcode_type, 16#07#),
      2249 => to_slv(opcode_type, 16#06#),
      2250 => to_slv(opcode_type, 16#02#),
      2251 => to_slv(opcode_type, 16#0B#),
      2252 => to_slv(opcode_type, 16#07#),
      2253 => to_slv(opcode_type, 16#0F#),
      2254 => to_slv(opcode_type, 16#0D#),
      2255 => to_slv(opcode_type, 16#06#),
      2256 => to_slv(opcode_type, 16#09#),
      2257 => to_slv(opcode_type, 16#10#),
      2258 => to_slv(opcode_type, 16#0C#),
      2259 => to_slv(opcode_type, 16#09#),
      2260 => to_slv(opcode_type, 16#0F#),
      2261 => to_slv(opcode_type, 16#D6#),
      2262 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#08#),
      2273 => to_slv(opcode_type, 16#09#),
      2274 => to_slv(opcode_type, 16#01#),
      2275 => to_slv(opcode_type, 16#05#),
      2276 => to_slv(opcode_type, 16#0C#),
      2277 => to_slv(opcode_type, 16#08#),
      2278 => to_slv(opcode_type, 16#08#),
      2279 => to_slv(opcode_type, 16#11#),
      2280 => to_slv(opcode_type, 16#0C#),
      2281 => to_slv(opcode_type, 16#04#),
      2282 => to_slv(opcode_type, 16#F8#),
      2283 => to_slv(opcode_type, 16#08#),
      2284 => to_slv(opcode_type, 16#03#),
      2285 => to_slv(opcode_type, 16#02#),
      2286 => to_slv(opcode_type, 16#0B#),
      2287 => to_slv(opcode_type, 16#09#),
      2288 => to_slv(opcode_type, 16#08#),
      2289 => to_slv(opcode_type, 16#0F#),
      2290 => to_slv(opcode_type, 16#11#),
      2291 => to_slv(opcode_type, 16#09#),
      2292 => to_slv(opcode_type, 16#11#),
      2293 => to_slv(opcode_type, 16#0E#),
      2294 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#07#),
      2305 => to_slv(opcode_type, 16#03#),
      2306 => to_slv(opcode_type, 16#06#),
      2307 => to_slv(opcode_type, 16#03#),
      2308 => to_slv(opcode_type, 16#11#),
      2309 => to_slv(opcode_type, 16#09#),
      2310 => to_slv(opcode_type, 16#0A#),
      2311 => to_slv(opcode_type, 16#0D#),
      2312 => to_slv(opcode_type, 16#08#),
      2313 => to_slv(opcode_type, 16#08#),
      2314 => to_slv(opcode_type, 16#09#),
      2315 => to_slv(opcode_type, 16#0D#),
      2316 => to_slv(opcode_type, 16#0C#),
      2317 => to_slv(opcode_type, 16#08#),
      2318 => to_slv(opcode_type, 16#0D#),
      2319 => to_slv(opcode_type, 16#B9#),
      2320 => to_slv(opcode_type, 16#07#),
      2321 => to_slv(opcode_type, 16#08#),
      2322 => to_slv(opcode_type, 16#0D#),
      2323 => to_slv(opcode_type, 16#0E#),
      2324 => to_slv(opcode_type, 16#04#),
      2325 => to_slv(opcode_type, 16#0E#),
      2326 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#09#),
      2337 => to_slv(opcode_type, 16#04#),
      2338 => to_slv(opcode_type, 16#08#),
      2339 => to_slv(opcode_type, 16#01#),
      2340 => to_slv(opcode_type, 16#0C#),
      2341 => to_slv(opcode_type, 16#03#),
      2342 => to_slv(opcode_type, 16#10#),
      2343 => to_slv(opcode_type, 16#07#),
      2344 => to_slv(opcode_type, 16#08#),
      2345 => to_slv(opcode_type, 16#08#),
      2346 => to_slv(opcode_type, 16#0C#),
      2347 => to_slv(opcode_type, 16#10#),
      2348 => to_slv(opcode_type, 16#07#),
      2349 => to_slv(opcode_type, 16#0C#),
      2350 => to_slv(opcode_type, 16#10#),
      2351 => to_slv(opcode_type, 16#08#),
      2352 => to_slv(opcode_type, 16#08#),
      2353 => to_slv(opcode_type, 16#1F#),
      2354 => to_slv(opcode_type, 16#0D#),
      2355 => to_slv(opcode_type, 16#07#),
      2356 => to_slv(opcode_type, 16#0E#),
      2357 => to_slv(opcode_type, 16#11#),
      2358 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#08#),
      2369 => to_slv(opcode_type, 16#06#),
      2370 => to_slv(opcode_type, 16#08#),
      2371 => to_slv(opcode_type, 16#07#),
      2372 => to_slv(opcode_type, 16#0D#),
      2373 => to_slv(opcode_type, 16#0F#),
      2374 => to_slv(opcode_type, 16#05#),
      2375 => to_slv(opcode_type, 16#0F#),
      2376 => to_slv(opcode_type, 16#02#),
      2377 => to_slv(opcode_type, 16#09#),
      2378 => to_slv(opcode_type, 16#10#),
      2379 => to_slv(opcode_type, 16#0E#),
      2380 => to_slv(opcode_type, 16#09#),
      2381 => to_slv(opcode_type, 16#07#),
      2382 => to_slv(opcode_type, 16#03#),
      2383 => to_slv(opcode_type, 16#0D#),
      2384 => to_slv(opcode_type, 16#04#),
      2385 => to_slv(opcode_type, 16#0F#),
      2386 => to_slv(opcode_type, 16#04#),
      2387 => to_slv(opcode_type, 16#08#),
      2388 => to_slv(opcode_type, 16#0B#),
      2389 => to_slv(opcode_type, 16#7A#),
      2390 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#08#),
      2401 => to_slv(opcode_type, 16#09#),
      2402 => to_slv(opcode_type, 16#05#),
      2403 => to_slv(opcode_type, 16#05#),
      2404 => to_slv(opcode_type, 16#11#),
      2405 => to_slv(opcode_type, 16#03#),
      2406 => to_slv(opcode_type, 16#06#),
      2407 => to_slv(opcode_type, 16#0E#),
      2408 => to_slv(opcode_type, 16#0A#),
      2409 => to_slv(opcode_type, 16#06#),
      2410 => to_slv(opcode_type, 16#07#),
      2411 => to_slv(opcode_type, 16#09#),
      2412 => to_slv(opcode_type, 16#0C#),
      2413 => to_slv(opcode_type, 16#0B#),
      2414 => to_slv(opcode_type, 16#04#),
      2415 => to_slv(opcode_type, 16#11#),
      2416 => to_slv(opcode_type, 16#07#),
      2417 => to_slv(opcode_type, 16#08#),
      2418 => to_slv(opcode_type, 16#C6#),
      2419 => to_slv(opcode_type, 16#0F#),
      2420 => to_slv(opcode_type, 16#02#),
      2421 => to_slv(opcode_type, 16#0D#),
      2422 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#08#),
      2433 => to_slv(opcode_type, 16#07#),
      2434 => to_slv(opcode_type, 16#03#),
      2435 => to_slv(opcode_type, 16#03#),
      2436 => to_slv(opcode_type, 16#11#),
      2437 => to_slv(opcode_type, 16#03#),
      2438 => to_slv(opcode_type, 16#01#),
      2439 => to_slv(opcode_type, 16#0A#),
      2440 => to_slv(opcode_type, 16#07#),
      2441 => to_slv(opcode_type, 16#06#),
      2442 => to_slv(opcode_type, 16#04#),
      2443 => to_slv(opcode_type, 16#0F#),
      2444 => to_slv(opcode_type, 16#07#),
      2445 => to_slv(opcode_type, 16#11#),
      2446 => to_slv(opcode_type, 16#0D#),
      2447 => to_slv(opcode_type, 16#07#),
      2448 => to_slv(opcode_type, 16#08#),
      2449 => to_slv(opcode_type, 16#0A#),
      2450 => to_slv(opcode_type, 16#0B#),
      2451 => to_slv(opcode_type, 16#07#),
      2452 => to_slv(opcode_type, 16#0E#),
      2453 => to_slv(opcode_type, 16#11#),
      2454 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#09#),
      2465 => to_slv(opcode_type, 16#04#),
      2466 => to_slv(opcode_type, 16#09#),
      2467 => to_slv(opcode_type, 16#06#),
      2468 => to_slv(opcode_type, 16#2F#),
      2469 => to_slv(opcode_type, 16#11#),
      2470 => to_slv(opcode_type, 16#07#),
      2471 => to_slv(opcode_type, 16#5A#),
      2472 => to_slv(opcode_type, 16#0C#),
      2473 => to_slv(opcode_type, 16#09#),
      2474 => to_slv(opcode_type, 16#07#),
      2475 => to_slv(opcode_type, 16#02#),
      2476 => to_slv(opcode_type, 16#0F#),
      2477 => to_slv(opcode_type, 16#05#),
      2478 => to_slv(opcode_type, 16#0C#),
      2479 => to_slv(opcode_type, 16#07#),
      2480 => to_slv(opcode_type, 16#07#),
      2481 => to_slv(opcode_type, 16#0E#),
      2482 => to_slv(opcode_type, 16#0D#),
      2483 => to_slv(opcode_type, 16#07#),
      2484 => to_slv(opcode_type, 16#0E#),
      2485 => to_slv(opcode_type, 16#0A#),
      2486 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#06#),
      2497 => to_slv(opcode_type, 16#08#),
      2498 => to_slv(opcode_type, 16#04#),
      2499 => to_slv(opcode_type, 16#06#),
      2500 => to_slv(opcode_type, 16#11#),
      2501 => to_slv(opcode_type, 16#CE#),
      2502 => to_slv(opcode_type, 16#09#),
      2503 => to_slv(opcode_type, 16#04#),
      2504 => to_slv(opcode_type, 16#0A#),
      2505 => to_slv(opcode_type, 16#06#),
      2506 => to_slv(opcode_type, 16#11#),
      2507 => to_slv(opcode_type, 16#0C#),
      2508 => to_slv(opcode_type, 16#06#),
      2509 => to_slv(opcode_type, 16#04#),
      2510 => to_slv(opcode_type, 16#09#),
      2511 => to_slv(opcode_type, 16#0B#),
      2512 => to_slv(opcode_type, 16#0A#),
      2513 => to_slv(opcode_type, 16#07#),
      2514 => to_slv(opcode_type, 16#06#),
      2515 => to_slv(opcode_type, 16#0C#),
      2516 => to_slv(opcode_type, 16#0A#),
      2517 => to_slv(opcode_type, 16#0D#),
      2518 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#02#),
      2530 => to_slv(opcode_type, 16#07#),
      2531 => to_slv(opcode_type, 16#08#),
      2532 => to_slv(opcode_type, 16#11#),
      2533 => to_slv(opcode_type, 16#0A#),
      2534 => to_slv(opcode_type, 16#09#),
      2535 => to_slv(opcode_type, 16#11#),
      2536 => to_slv(opcode_type, 16#0C#),
      2537 => to_slv(opcode_type, 16#08#),
      2538 => to_slv(opcode_type, 16#08#),
      2539 => to_slv(opcode_type, 16#06#),
      2540 => to_slv(opcode_type, 16#10#),
      2541 => to_slv(opcode_type, 16#6C#),
      2542 => to_slv(opcode_type, 16#06#),
      2543 => to_slv(opcode_type, 16#11#),
      2544 => to_slv(opcode_type, 16#0E#),
      2545 => to_slv(opcode_type, 16#09#),
      2546 => to_slv(opcode_type, 16#03#),
      2547 => to_slv(opcode_type, 16#10#),
      2548 => to_slv(opcode_type, 16#03#),
      2549 => to_slv(opcode_type, 16#0E#),
      2550 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#06#),
      2561 => to_slv(opcode_type, 16#01#),
      2562 => to_slv(opcode_type, 16#06#),
      2563 => to_slv(opcode_type, 16#08#),
      2564 => to_slv(opcode_type, 16#0D#),
      2565 => to_slv(opcode_type, 16#0B#),
      2566 => to_slv(opcode_type, 16#08#),
      2567 => to_slv(opcode_type, 16#0C#),
      2568 => to_slv(opcode_type, 16#10#),
      2569 => to_slv(opcode_type, 16#09#),
      2570 => to_slv(opcode_type, 16#08#),
      2571 => to_slv(opcode_type, 16#07#),
      2572 => to_slv(opcode_type, 16#0B#),
      2573 => to_slv(opcode_type, 16#10#),
      2574 => to_slv(opcode_type, 16#01#),
      2575 => to_slv(opcode_type, 16#0B#),
      2576 => to_slv(opcode_type, 16#08#),
      2577 => to_slv(opcode_type, 16#04#),
      2578 => to_slv(opcode_type, 16#0F#),
      2579 => to_slv(opcode_type, 16#08#),
      2580 => to_slv(opcode_type, 16#0E#),
      2581 => to_slv(opcode_type, 16#0C#),
      2582 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#06#),
      2593 => to_slv(opcode_type, 16#09#),
      2594 => to_slv(opcode_type, 16#07#),
      2595 => to_slv(opcode_type, 16#04#),
      2596 => to_slv(opcode_type, 16#0B#),
      2597 => to_slv(opcode_type, 16#08#),
      2598 => to_slv(opcode_type, 16#10#),
      2599 => to_slv(opcode_type, 16#11#),
      2600 => to_slv(opcode_type, 16#09#),
      2601 => to_slv(opcode_type, 16#02#),
      2602 => to_slv(opcode_type, 16#10#),
      2603 => to_slv(opcode_type, 16#07#),
      2604 => to_slv(opcode_type, 16#0F#),
      2605 => to_slv(opcode_type, 16#11#),
      2606 => to_slv(opcode_type, 16#04#),
      2607 => to_slv(opcode_type, 16#06#),
      2608 => to_slv(opcode_type, 16#06#),
      2609 => to_slv(opcode_type, 16#0B#),
      2610 => to_slv(opcode_type, 16#11#),
      2611 => to_slv(opcode_type, 16#07#),
      2612 => to_slv(opcode_type, 16#11#),
      2613 => to_slv(opcode_type, 16#0C#),
      2614 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#08#),
      2625 => to_slv(opcode_type, 16#06#),
      2626 => to_slv(opcode_type, 16#08#),
      2627 => to_slv(opcode_type, 16#02#),
      2628 => to_slv(opcode_type, 16#0D#),
      2629 => to_slv(opcode_type, 16#01#),
      2630 => to_slv(opcode_type, 16#E0#),
      2631 => to_slv(opcode_type, 16#03#),
      2632 => to_slv(opcode_type, 16#07#),
      2633 => to_slv(opcode_type, 16#10#),
      2634 => to_slv(opcode_type, 16#0B#),
      2635 => to_slv(opcode_type, 16#07#),
      2636 => to_slv(opcode_type, 16#01#),
      2637 => to_slv(opcode_type, 16#02#),
      2638 => to_slv(opcode_type, 16#10#),
      2639 => to_slv(opcode_type, 16#06#),
      2640 => to_slv(opcode_type, 16#06#),
      2641 => to_slv(opcode_type, 16#0C#),
      2642 => to_slv(opcode_type, 16#0D#),
      2643 => to_slv(opcode_type, 16#09#),
      2644 => to_slv(opcode_type, 16#0C#),
      2645 => to_slv(opcode_type, 16#0C#),
      2646 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#09#),
      2657 => to_slv(opcode_type, 16#01#),
      2658 => to_slv(opcode_type, 16#09#),
      2659 => to_slv(opcode_type, 16#07#),
      2660 => to_slv(opcode_type, 16#0C#),
      2661 => to_slv(opcode_type, 16#11#),
      2662 => to_slv(opcode_type, 16#02#),
      2663 => to_slv(opcode_type, 16#0D#),
      2664 => to_slv(opcode_type, 16#06#),
      2665 => to_slv(opcode_type, 16#07#),
      2666 => to_slv(opcode_type, 16#06#),
      2667 => to_slv(opcode_type, 16#0B#),
      2668 => to_slv(opcode_type, 16#84#),
      2669 => to_slv(opcode_type, 16#02#),
      2670 => to_slv(opcode_type, 16#0D#),
      2671 => to_slv(opcode_type, 16#06#),
      2672 => to_slv(opcode_type, 16#08#),
      2673 => to_slv(opcode_type, 16#0D#),
      2674 => to_slv(opcode_type, 16#10#),
      2675 => to_slv(opcode_type, 16#09#),
      2676 => to_slv(opcode_type, 16#0B#),
      2677 => to_slv(opcode_type, 16#0B#),
      2678 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#09#),
      2689 => to_slv(opcode_type, 16#09#),
      2690 => to_slv(opcode_type, 16#08#),
      2691 => to_slv(opcode_type, 16#08#),
      2692 => to_slv(opcode_type, 16#0E#),
      2693 => to_slv(opcode_type, 16#0D#),
      2694 => to_slv(opcode_type, 16#03#),
      2695 => to_slv(opcode_type, 16#0B#),
      2696 => to_slv(opcode_type, 16#06#),
      2697 => to_slv(opcode_type, 16#07#),
      2698 => to_slv(opcode_type, 16#11#),
      2699 => to_slv(opcode_type, 16#0A#),
      2700 => to_slv(opcode_type, 16#04#),
      2701 => to_slv(opcode_type, 16#ED#),
      2702 => to_slv(opcode_type, 16#01#),
      2703 => to_slv(opcode_type, 16#07#),
      2704 => to_slv(opcode_type, 16#08#),
      2705 => to_slv(opcode_type, 16#0C#),
      2706 => to_slv(opcode_type, 16#0C#),
      2707 => to_slv(opcode_type, 16#06#),
      2708 => to_slv(opcode_type, 16#0A#),
      2709 => to_slv(opcode_type, 16#0C#),
      2710 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#08#),
      2721 => to_slv(opcode_type, 16#03#),
      2722 => to_slv(opcode_type, 16#06#),
      2723 => to_slv(opcode_type, 16#01#),
      2724 => to_slv(opcode_type, 16#10#),
      2725 => to_slv(opcode_type, 16#07#),
      2726 => to_slv(opcode_type, 16#0D#),
      2727 => to_slv(opcode_type, 16#0A#),
      2728 => to_slv(opcode_type, 16#07#),
      2729 => to_slv(opcode_type, 16#06#),
      2730 => to_slv(opcode_type, 16#01#),
      2731 => to_slv(opcode_type, 16#0F#),
      2732 => to_slv(opcode_type, 16#07#),
      2733 => to_slv(opcode_type, 16#10#),
      2734 => to_slv(opcode_type, 16#0B#),
      2735 => to_slv(opcode_type, 16#07#),
      2736 => to_slv(opcode_type, 16#08#),
      2737 => to_slv(opcode_type, 16#0F#),
      2738 => to_slv(opcode_type, 16#0F#),
      2739 => to_slv(opcode_type, 16#06#),
      2740 => to_slv(opcode_type, 16#0D#),
      2741 => to_slv(opcode_type, 16#0A#),
      2742 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#06#),
      2753 => to_slv(opcode_type, 16#02#),
      2754 => to_slv(opcode_type, 16#08#),
      2755 => to_slv(opcode_type, 16#05#),
      2756 => to_slv(opcode_type, 16#11#),
      2757 => to_slv(opcode_type, 16#03#),
      2758 => to_slv(opcode_type, 16#0A#),
      2759 => to_slv(opcode_type, 16#06#),
      2760 => to_slv(opcode_type, 16#06#),
      2761 => to_slv(opcode_type, 16#08#),
      2762 => to_slv(opcode_type, 16#0F#),
      2763 => to_slv(opcode_type, 16#0A#),
      2764 => to_slv(opcode_type, 16#06#),
      2765 => to_slv(opcode_type, 16#0F#),
      2766 => to_slv(opcode_type, 16#F5#),
      2767 => to_slv(opcode_type, 16#06#),
      2768 => to_slv(opcode_type, 16#06#),
      2769 => to_slv(opcode_type, 16#0B#),
      2770 => to_slv(opcode_type, 16#0D#),
      2771 => to_slv(opcode_type, 16#09#),
      2772 => to_slv(opcode_type, 16#11#),
      2773 => to_slv(opcode_type, 16#0F#),
      2774 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#09#),
      2785 => to_slv(opcode_type, 16#02#),
      2786 => to_slv(opcode_type, 16#09#),
      2787 => to_slv(opcode_type, 16#06#),
      2788 => to_slv(opcode_type, 16#0E#),
      2789 => to_slv(opcode_type, 16#1B#),
      2790 => to_slv(opcode_type, 16#06#),
      2791 => to_slv(opcode_type, 16#11#),
      2792 => to_slv(opcode_type, 16#C2#),
      2793 => to_slv(opcode_type, 16#06#),
      2794 => to_slv(opcode_type, 16#06#),
      2795 => to_slv(opcode_type, 16#08#),
      2796 => to_slv(opcode_type, 16#0B#),
      2797 => to_slv(opcode_type, 16#11#),
      2798 => to_slv(opcode_type, 16#06#),
      2799 => to_slv(opcode_type, 16#10#),
      2800 => to_slv(opcode_type, 16#0F#),
      2801 => to_slv(opcode_type, 16#07#),
      2802 => to_slv(opcode_type, 16#04#),
      2803 => to_slv(opcode_type, 16#0D#),
      2804 => to_slv(opcode_type, 16#03#),
      2805 => to_slv(opcode_type, 16#0F#),
      2806 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#06#),
      2817 => to_slv(opcode_type, 16#07#),
      2818 => to_slv(opcode_type, 16#07#),
      2819 => to_slv(opcode_type, 16#06#),
      2820 => to_slv(opcode_type, 16#11#),
      2821 => to_slv(opcode_type, 16#6E#),
      2822 => to_slv(opcode_type, 16#05#),
      2823 => to_slv(opcode_type, 16#11#),
      2824 => to_slv(opcode_type, 16#08#),
      2825 => to_slv(opcode_type, 16#05#),
      2826 => to_slv(opcode_type, 16#0B#),
      2827 => to_slv(opcode_type, 16#01#),
      2828 => to_slv(opcode_type, 16#0C#),
      2829 => to_slv(opcode_type, 16#09#),
      2830 => to_slv(opcode_type, 16#05#),
      2831 => to_slv(opcode_type, 16#02#),
      2832 => to_slv(opcode_type, 16#0F#),
      2833 => to_slv(opcode_type, 16#06#),
      2834 => to_slv(opcode_type, 16#08#),
      2835 => to_slv(opcode_type, 16#11#),
      2836 => to_slv(opcode_type, 16#0E#),
      2837 => to_slv(opcode_type, 16#0B#),
      2838 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#06#),
      2849 => to_slv(opcode_type, 16#03#),
      2850 => to_slv(opcode_type, 16#06#),
      2851 => to_slv(opcode_type, 16#08#),
      2852 => to_slv(opcode_type, 16#11#),
      2853 => to_slv(opcode_type, 16#0E#),
      2854 => to_slv(opcode_type, 16#05#),
      2855 => to_slv(opcode_type, 16#0B#),
      2856 => to_slv(opcode_type, 16#07#),
      2857 => to_slv(opcode_type, 16#08#),
      2858 => to_slv(opcode_type, 16#05#),
      2859 => to_slv(opcode_type, 16#10#),
      2860 => to_slv(opcode_type, 16#06#),
      2861 => to_slv(opcode_type, 16#10#),
      2862 => to_slv(opcode_type, 16#0F#),
      2863 => to_slv(opcode_type, 16#07#),
      2864 => to_slv(opcode_type, 16#06#),
      2865 => to_slv(opcode_type, 16#0C#),
      2866 => to_slv(opcode_type, 16#0C#),
      2867 => to_slv(opcode_type, 16#07#),
      2868 => to_slv(opcode_type, 16#0D#),
      2869 => to_slv(opcode_type, 16#11#),
      2870 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#07#),
      2881 => to_slv(opcode_type, 16#06#),
      2882 => to_slv(opcode_type, 16#06#),
      2883 => to_slv(opcode_type, 16#08#),
      2884 => to_slv(opcode_type, 16#10#),
      2885 => to_slv(opcode_type, 16#0F#),
      2886 => to_slv(opcode_type, 16#08#),
      2887 => to_slv(opcode_type, 16#10#),
      2888 => to_slv(opcode_type, 16#0D#),
      2889 => to_slv(opcode_type, 16#04#),
      2890 => to_slv(opcode_type, 16#06#),
      2891 => to_slv(opcode_type, 16#0E#),
      2892 => to_slv(opcode_type, 16#10#),
      2893 => to_slv(opcode_type, 16#06#),
      2894 => to_slv(opcode_type, 16#09#),
      2895 => to_slv(opcode_type, 16#05#),
      2896 => to_slv(opcode_type, 16#0B#),
      2897 => to_slv(opcode_type, 16#09#),
      2898 => to_slv(opcode_type, 16#0C#),
      2899 => to_slv(opcode_type, 16#0F#),
      2900 => to_slv(opcode_type, 16#01#),
      2901 => to_slv(opcode_type, 16#0E#),
      2902 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#06#),
      2913 => to_slv(opcode_type, 16#07#),
      2914 => to_slv(opcode_type, 16#04#),
      2915 => to_slv(opcode_type, 16#09#),
      2916 => to_slv(opcode_type, 16#0C#),
      2917 => to_slv(opcode_type, 16#0D#),
      2918 => to_slv(opcode_type, 16#08#),
      2919 => to_slv(opcode_type, 16#02#),
      2920 => to_slv(opcode_type, 16#0F#),
      2921 => to_slv(opcode_type, 16#07#),
      2922 => to_slv(opcode_type, 16#B1#),
      2923 => to_slv(opcode_type, 16#11#),
      2924 => to_slv(opcode_type, 16#09#),
      2925 => to_slv(opcode_type, 16#02#),
      2926 => to_slv(opcode_type, 16#08#),
      2927 => to_slv(opcode_type, 16#0C#),
      2928 => to_slv(opcode_type, 16#0E#),
      2929 => to_slv(opcode_type, 16#07#),
      2930 => to_slv(opcode_type, 16#08#),
      2931 => to_slv(opcode_type, 16#0C#),
      2932 => to_slv(opcode_type, 16#0F#),
      2933 => to_slv(opcode_type, 16#0E#),
      2934 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#08#),
      2945 => to_slv(opcode_type, 16#07#),
      2946 => to_slv(opcode_type, 16#03#),
      2947 => to_slv(opcode_type, 16#03#),
      2948 => to_slv(opcode_type, 16#0D#),
      2949 => to_slv(opcode_type, 16#09#),
      2950 => to_slv(opcode_type, 16#09#),
      2951 => to_slv(opcode_type, 16#12#),
      2952 => to_slv(opcode_type, 16#11#),
      2953 => to_slv(opcode_type, 16#08#),
      2954 => to_slv(opcode_type, 16#10#),
      2955 => to_slv(opcode_type, 16#0E#),
      2956 => to_slv(opcode_type, 16#08#),
      2957 => to_slv(opcode_type, 16#02#),
      2958 => to_slv(opcode_type, 16#05#),
      2959 => to_slv(opcode_type, 16#0A#),
      2960 => to_slv(opcode_type, 16#08#),
      2961 => to_slv(opcode_type, 16#02#),
      2962 => to_slv(opcode_type, 16#10#),
      2963 => to_slv(opcode_type, 16#09#),
      2964 => to_slv(opcode_type, 16#0C#),
      2965 => to_slv(opcode_type, 16#0E#),
      2966 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#08#),
      2977 => to_slv(opcode_type, 16#02#),
      2978 => to_slv(opcode_type, 16#06#),
      2979 => to_slv(opcode_type, 16#05#),
      2980 => to_slv(opcode_type, 16#10#),
      2981 => to_slv(opcode_type, 16#03#),
      2982 => to_slv(opcode_type, 16#DB#),
      2983 => to_slv(opcode_type, 16#08#),
      2984 => to_slv(opcode_type, 16#06#),
      2985 => to_slv(opcode_type, 16#06#),
      2986 => to_slv(opcode_type, 16#11#),
      2987 => to_slv(opcode_type, 16#0C#),
      2988 => to_slv(opcode_type, 16#07#),
      2989 => to_slv(opcode_type, 16#0D#),
      2990 => to_slv(opcode_type, 16#45#),
      2991 => to_slv(opcode_type, 16#09#),
      2992 => to_slv(opcode_type, 16#07#),
      2993 => to_slv(opcode_type, 16#0F#),
      2994 => to_slv(opcode_type, 16#11#),
      2995 => to_slv(opcode_type, 16#09#),
      2996 => to_slv(opcode_type, 16#0A#),
      2997 => to_slv(opcode_type, 16#0D#),
      2998 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#06#),
      3009 => to_slv(opcode_type, 16#08#),
      3010 => to_slv(opcode_type, 16#02#),
      3011 => to_slv(opcode_type, 16#02#),
      3012 => to_slv(opcode_type, 16#0D#),
      3013 => to_slv(opcode_type, 16#01#),
      3014 => to_slv(opcode_type, 16#09#),
      3015 => to_slv(opcode_type, 16#0C#),
      3016 => to_slv(opcode_type, 16#0C#),
      3017 => to_slv(opcode_type, 16#06#),
      3018 => to_slv(opcode_type, 16#06#),
      3019 => to_slv(opcode_type, 16#06#),
      3020 => to_slv(opcode_type, 16#10#),
      3021 => to_slv(opcode_type, 16#0B#),
      3022 => to_slv(opcode_type, 16#07#),
      3023 => to_slv(opcode_type, 16#0E#),
      3024 => to_slv(opcode_type, 16#7C#),
      3025 => to_slv(opcode_type, 16#06#),
      3026 => to_slv(opcode_type, 16#01#),
      3027 => to_slv(opcode_type, 16#61#),
      3028 => to_slv(opcode_type, 16#05#),
      3029 => to_slv(opcode_type, 16#0B#),
      3030 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#08#),
      3041 => to_slv(opcode_type, 16#05#),
      3042 => to_slv(opcode_type, 16#07#),
      3043 => to_slv(opcode_type, 16#05#),
      3044 => to_slv(opcode_type, 16#10#),
      3045 => to_slv(opcode_type, 16#01#),
      3046 => to_slv(opcode_type, 16#0C#),
      3047 => to_slv(opcode_type, 16#09#),
      3048 => to_slv(opcode_type, 16#08#),
      3049 => to_slv(opcode_type, 16#06#),
      3050 => to_slv(opcode_type, 16#10#),
      3051 => to_slv(opcode_type, 16#0A#),
      3052 => to_slv(opcode_type, 16#09#),
      3053 => to_slv(opcode_type, 16#0E#),
      3054 => to_slv(opcode_type, 16#0A#),
      3055 => to_slv(opcode_type, 16#08#),
      3056 => to_slv(opcode_type, 16#06#),
      3057 => to_slv(opcode_type, 16#0F#),
      3058 => to_slv(opcode_type, 16#10#),
      3059 => to_slv(opcode_type, 16#09#),
      3060 => to_slv(opcode_type, 16#0C#),
      3061 => to_slv(opcode_type, 16#11#),
      3062 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#06#),
      3073 => to_slv(opcode_type, 16#04#),
      3074 => to_slv(opcode_type, 16#06#),
      3075 => to_slv(opcode_type, 16#02#),
      3076 => to_slv(opcode_type, 16#0A#),
      3077 => to_slv(opcode_type, 16#02#),
      3078 => to_slv(opcode_type, 16#0E#),
      3079 => to_slv(opcode_type, 16#08#),
      3080 => to_slv(opcode_type, 16#09#),
      3081 => to_slv(opcode_type, 16#07#),
      3082 => to_slv(opcode_type, 16#10#),
      3083 => to_slv(opcode_type, 16#11#),
      3084 => to_slv(opcode_type, 16#08#),
      3085 => to_slv(opcode_type, 16#0D#),
      3086 => to_slv(opcode_type, 16#74#),
      3087 => to_slv(opcode_type, 16#08#),
      3088 => to_slv(opcode_type, 16#07#),
      3089 => to_slv(opcode_type, 16#0E#),
      3090 => to_slv(opcode_type, 16#10#),
      3091 => to_slv(opcode_type, 16#06#),
      3092 => to_slv(opcode_type, 16#11#),
      3093 => to_slv(opcode_type, 16#10#),
      3094 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#07#),
      3105 => to_slv(opcode_type, 16#01#),
      3106 => to_slv(opcode_type, 16#08#),
      3107 => to_slv(opcode_type, 16#07#),
      3108 => to_slv(opcode_type, 16#0D#),
      3109 => to_slv(opcode_type, 16#0B#),
      3110 => to_slv(opcode_type, 16#09#),
      3111 => to_slv(opcode_type, 16#0D#),
      3112 => to_slv(opcode_type, 16#AC#),
      3113 => to_slv(opcode_type, 16#08#),
      3114 => to_slv(opcode_type, 16#08#),
      3115 => to_slv(opcode_type, 16#01#),
      3116 => to_slv(opcode_type, 16#10#),
      3117 => to_slv(opcode_type, 16#06#),
      3118 => to_slv(opcode_type, 16#0E#),
      3119 => to_slv(opcode_type, 16#10#),
      3120 => to_slv(opcode_type, 16#07#),
      3121 => to_slv(opcode_type, 16#05#),
      3122 => to_slv(opcode_type, 16#0B#),
      3123 => to_slv(opcode_type, 16#07#),
      3124 => to_slv(opcode_type, 16#0A#),
      3125 => to_slv(opcode_type, 16#10#),
      3126 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#07#),
      3137 => to_slv(opcode_type, 16#02#),
      3138 => to_slv(opcode_type, 16#07#),
      3139 => to_slv(opcode_type, 16#01#),
      3140 => to_slv(opcode_type, 16#0C#),
      3141 => to_slv(opcode_type, 16#06#),
      3142 => to_slv(opcode_type, 16#0D#),
      3143 => to_slv(opcode_type, 16#11#),
      3144 => to_slv(opcode_type, 16#08#),
      3145 => to_slv(opcode_type, 16#09#),
      3146 => to_slv(opcode_type, 16#05#),
      3147 => to_slv(opcode_type, 16#0D#),
      3148 => to_slv(opcode_type, 16#06#),
      3149 => to_slv(opcode_type, 16#0F#),
      3150 => to_slv(opcode_type, 16#0F#),
      3151 => to_slv(opcode_type, 16#09#),
      3152 => to_slv(opcode_type, 16#08#),
      3153 => to_slv(opcode_type, 16#0E#),
      3154 => to_slv(opcode_type, 16#0E#),
      3155 => to_slv(opcode_type, 16#08#),
      3156 => to_slv(opcode_type, 16#0A#),
      3157 => to_slv(opcode_type, 16#11#),
      3158 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#09#),
      3169 => to_slv(opcode_type, 16#08#),
      3170 => to_slv(opcode_type, 16#03#),
      3171 => to_slv(opcode_type, 16#05#),
      3172 => to_slv(opcode_type, 16#11#),
      3173 => to_slv(opcode_type, 16#02#),
      3174 => to_slv(opcode_type, 16#03#),
      3175 => to_slv(opcode_type, 16#0F#),
      3176 => to_slv(opcode_type, 16#07#),
      3177 => to_slv(opcode_type, 16#08#),
      3178 => to_slv(opcode_type, 16#07#),
      3179 => to_slv(opcode_type, 16#0D#),
      3180 => to_slv(opcode_type, 16#0E#),
      3181 => to_slv(opcode_type, 16#03#),
      3182 => to_slv(opcode_type, 16#10#),
      3183 => to_slv(opcode_type, 16#06#),
      3184 => to_slv(opcode_type, 16#09#),
      3185 => to_slv(opcode_type, 16#0F#),
      3186 => to_slv(opcode_type, 16#73#),
      3187 => to_slv(opcode_type, 16#07#),
      3188 => to_slv(opcode_type, 16#0F#),
      3189 => to_slv(opcode_type, 16#0D#),
      3190 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#06#),
      3201 => to_slv(opcode_type, 16#02#),
      3202 => to_slv(opcode_type, 16#06#),
      3203 => to_slv(opcode_type, 16#05#),
      3204 => to_slv(opcode_type, 16#99#),
      3205 => to_slv(opcode_type, 16#06#),
      3206 => to_slv(opcode_type, 16#A1#),
      3207 => to_slv(opcode_type, 16#0C#),
      3208 => to_slv(opcode_type, 16#08#),
      3209 => to_slv(opcode_type, 16#09#),
      3210 => to_slv(opcode_type, 16#03#),
      3211 => to_slv(opcode_type, 16#10#),
      3212 => to_slv(opcode_type, 16#06#),
      3213 => to_slv(opcode_type, 16#0D#),
      3214 => to_slv(opcode_type, 16#0B#),
      3215 => to_slv(opcode_type, 16#06#),
      3216 => to_slv(opcode_type, 16#08#),
      3217 => to_slv(opcode_type, 16#10#),
      3218 => to_slv(opcode_type, 16#0A#),
      3219 => to_slv(opcode_type, 16#08#),
      3220 => to_slv(opcode_type, 16#0E#),
      3221 => to_slv(opcode_type, 16#1B#),
      3222 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#08#),
      3233 => to_slv(opcode_type, 16#04#),
      3234 => to_slv(opcode_type, 16#06#),
      3235 => to_slv(opcode_type, 16#04#),
      3236 => to_slv(opcode_type, 16#0A#),
      3237 => to_slv(opcode_type, 16#09#),
      3238 => to_slv(opcode_type, 16#0A#),
      3239 => to_slv(opcode_type, 16#0A#),
      3240 => to_slv(opcode_type, 16#09#),
      3241 => to_slv(opcode_type, 16#07#),
      3242 => to_slv(opcode_type, 16#08#),
      3243 => to_slv(opcode_type, 16#0F#),
      3244 => to_slv(opcode_type, 16#0D#),
      3245 => to_slv(opcode_type, 16#09#),
      3246 => to_slv(opcode_type, 16#0B#),
      3247 => to_slv(opcode_type, 16#0A#),
      3248 => to_slv(opcode_type, 16#06#),
      3249 => to_slv(opcode_type, 16#03#),
      3250 => to_slv(opcode_type, 16#0F#),
      3251 => to_slv(opcode_type, 16#08#),
      3252 => to_slv(opcode_type, 16#0C#),
      3253 => to_slv(opcode_type, 16#0B#),
      3254 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#06#),
      3265 => to_slv(opcode_type, 16#06#),
      3266 => to_slv(opcode_type, 16#07#),
      3267 => to_slv(opcode_type, 16#01#),
      3268 => to_slv(opcode_type, 16#0D#),
      3269 => to_slv(opcode_type, 16#07#),
      3270 => to_slv(opcode_type, 16#10#),
      3271 => to_slv(opcode_type, 16#0B#),
      3272 => to_slv(opcode_type, 16#07#),
      3273 => to_slv(opcode_type, 16#03#),
      3274 => to_slv(opcode_type, 16#A8#),
      3275 => to_slv(opcode_type, 16#05#),
      3276 => to_slv(opcode_type, 16#0F#),
      3277 => to_slv(opcode_type, 16#08#),
      3278 => to_slv(opcode_type, 16#04#),
      3279 => to_slv(opcode_type, 16#07#),
      3280 => to_slv(opcode_type, 16#0D#),
      3281 => to_slv(opcode_type, 16#10#),
      3282 => to_slv(opcode_type, 16#02#),
      3283 => to_slv(opcode_type, 16#09#),
      3284 => to_slv(opcode_type, 16#0C#),
      3285 => to_slv(opcode_type, 16#11#),
      3286 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#06#),
      3297 => to_slv(opcode_type, 16#07#),
      3298 => to_slv(opcode_type, 16#09#),
      3299 => to_slv(opcode_type, 16#07#),
      3300 => to_slv(opcode_type, 16#10#),
      3301 => to_slv(opcode_type, 16#0F#),
      3302 => to_slv(opcode_type, 16#05#),
      3303 => to_slv(opcode_type, 16#0F#),
      3304 => to_slv(opcode_type, 16#06#),
      3305 => to_slv(opcode_type, 16#07#),
      3306 => to_slv(opcode_type, 16#11#),
      3307 => to_slv(opcode_type, 16#0B#),
      3308 => to_slv(opcode_type, 16#03#),
      3309 => to_slv(opcode_type, 16#0C#),
      3310 => to_slv(opcode_type, 16#05#),
      3311 => to_slv(opcode_type, 16#09#),
      3312 => to_slv(opcode_type, 16#06#),
      3313 => to_slv(opcode_type, 16#10#),
      3314 => to_slv(opcode_type, 16#0F#),
      3315 => to_slv(opcode_type, 16#06#),
      3316 => to_slv(opcode_type, 16#0B#),
      3317 => to_slv(opcode_type, 16#0D#),
      3318 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#07#),
      3329 => to_slv(opcode_type, 16#09#),
      3330 => to_slv(opcode_type, 16#03#),
      3331 => to_slv(opcode_type, 16#04#),
      3332 => to_slv(opcode_type, 16#0D#),
      3333 => to_slv(opcode_type, 16#09#),
      3334 => to_slv(opcode_type, 16#03#),
      3335 => to_slv(opcode_type, 16#0F#),
      3336 => to_slv(opcode_type, 16#05#),
      3337 => to_slv(opcode_type, 16#0C#),
      3338 => to_slv(opcode_type, 16#09#),
      3339 => to_slv(opcode_type, 16#06#),
      3340 => to_slv(opcode_type, 16#04#),
      3341 => to_slv(opcode_type, 16#0B#),
      3342 => to_slv(opcode_type, 16#01#),
      3343 => to_slv(opcode_type, 16#0C#),
      3344 => to_slv(opcode_type, 16#09#),
      3345 => to_slv(opcode_type, 16#08#),
      3346 => to_slv(opcode_type, 16#0A#),
      3347 => to_slv(opcode_type, 16#0F#),
      3348 => to_slv(opcode_type, 16#05#),
      3349 => to_slv(opcode_type, 16#10#),
      3350 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#08#),
      3361 => to_slv(opcode_type, 16#02#),
      3362 => to_slv(opcode_type, 16#07#),
      3363 => to_slv(opcode_type, 16#08#),
      3364 => to_slv(opcode_type, 16#10#),
      3365 => to_slv(opcode_type, 16#0E#),
      3366 => to_slv(opcode_type, 16#07#),
      3367 => to_slv(opcode_type, 16#7C#),
      3368 => to_slv(opcode_type, 16#0C#),
      3369 => to_slv(opcode_type, 16#07#),
      3370 => to_slv(opcode_type, 16#06#),
      3371 => to_slv(opcode_type, 16#01#),
      3372 => to_slv(opcode_type, 16#2B#),
      3373 => to_slv(opcode_type, 16#02#),
      3374 => to_slv(opcode_type, 16#0D#),
      3375 => to_slv(opcode_type, 16#08#),
      3376 => to_slv(opcode_type, 16#06#),
      3377 => to_slv(opcode_type, 16#A3#),
      3378 => to_slv(opcode_type, 16#0A#),
      3379 => to_slv(opcode_type, 16#06#),
      3380 => to_slv(opcode_type, 16#0F#),
      3381 => to_slv(opcode_type, 16#0B#),
      3382 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#09#),
      3393 => to_slv(opcode_type, 16#06#),
      3394 => to_slv(opcode_type, 16#08#),
      3395 => to_slv(opcode_type, 16#07#),
      3396 => to_slv(opcode_type, 16#11#),
      3397 => to_slv(opcode_type, 16#10#),
      3398 => to_slv(opcode_type, 16#07#),
      3399 => to_slv(opcode_type, 16#0A#),
      3400 => to_slv(opcode_type, 16#0F#),
      3401 => to_slv(opcode_type, 16#03#),
      3402 => to_slv(opcode_type, 16#06#),
      3403 => to_slv(opcode_type, 16#0B#),
      3404 => to_slv(opcode_type, 16#10#),
      3405 => to_slv(opcode_type, 16#06#),
      3406 => to_slv(opcode_type, 16#06#),
      3407 => to_slv(opcode_type, 16#08#),
      3408 => to_slv(opcode_type, 16#0F#),
      3409 => to_slv(opcode_type, 16#0B#),
      3410 => to_slv(opcode_type, 16#03#),
      3411 => to_slv(opcode_type, 16#0F#),
      3412 => to_slv(opcode_type, 16#02#),
      3413 => to_slv(opcode_type, 16#10#),
      3414 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#09#),
      3426 => to_slv(opcode_type, 16#09#),
      3427 => to_slv(opcode_type, 16#03#),
      3428 => to_slv(opcode_type, 16#0B#),
      3429 => to_slv(opcode_type, 16#05#),
      3430 => to_slv(opcode_type, 16#0A#),
      3431 => to_slv(opcode_type, 16#08#),
      3432 => to_slv(opcode_type, 16#07#),
      3433 => to_slv(opcode_type, 16#0C#),
      3434 => to_slv(opcode_type, 16#10#),
      3435 => to_slv(opcode_type, 16#08#),
      3436 => to_slv(opcode_type, 16#28#),
      3437 => to_slv(opcode_type, 16#95#),
      3438 => to_slv(opcode_type, 16#08#),
      3439 => to_slv(opcode_type, 16#03#),
      3440 => to_slv(opcode_type, 16#03#),
      3441 => to_slv(opcode_type, 16#0C#),
      3442 => to_slv(opcode_type, 16#04#),
      3443 => to_slv(opcode_type, 16#08#),
      3444 => to_slv(opcode_type, 16#0E#),
      3445 => to_slv(opcode_type, 16#0D#),
      3446 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#08#),
      3457 => to_slv(opcode_type, 16#03#),
      3458 => to_slv(opcode_type, 16#06#),
      3459 => to_slv(opcode_type, 16#07#),
      3460 => to_slv(opcode_type, 16#EE#),
      3461 => to_slv(opcode_type, 16#35#),
      3462 => to_slv(opcode_type, 16#03#),
      3463 => to_slv(opcode_type, 16#0A#),
      3464 => to_slv(opcode_type, 16#07#),
      3465 => to_slv(opcode_type, 16#09#),
      3466 => to_slv(opcode_type, 16#03#),
      3467 => to_slv(opcode_type, 16#0C#),
      3468 => to_slv(opcode_type, 16#06#),
      3469 => to_slv(opcode_type, 16#11#),
      3470 => to_slv(opcode_type, 16#0F#),
      3471 => to_slv(opcode_type, 16#09#),
      3472 => to_slv(opcode_type, 16#06#),
      3473 => to_slv(opcode_type, 16#0F#),
      3474 => to_slv(opcode_type, 16#0F#),
      3475 => to_slv(opcode_type, 16#08#),
      3476 => to_slv(opcode_type, 16#0C#),
      3477 => to_slv(opcode_type, 16#0F#),
      3478 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#09#),
      3489 => to_slv(opcode_type, 16#08#),
      3490 => to_slv(opcode_type, 16#05#),
      3491 => to_slv(opcode_type, 16#05#),
      3492 => to_slv(opcode_type, 16#0D#),
      3493 => to_slv(opcode_type, 16#04#),
      3494 => to_slv(opcode_type, 16#04#),
      3495 => to_slv(opcode_type, 16#0F#),
      3496 => to_slv(opcode_type, 16#08#),
      3497 => to_slv(opcode_type, 16#06#),
      3498 => to_slv(opcode_type, 16#05#),
      3499 => to_slv(opcode_type, 16#0A#),
      3500 => to_slv(opcode_type, 16#07#),
      3501 => to_slv(opcode_type, 16#0B#),
      3502 => to_slv(opcode_type, 16#11#),
      3503 => to_slv(opcode_type, 16#06#),
      3504 => to_slv(opcode_type, 16#09#),
      3505 => to_slv(opcode_type, 16#0E#),
      3506 => to_slv(opcode_type, 16#0E#),
      3507 => to_slv(opcode_type, 16#06#),
      3508 => to_slv(opcode_type, 16#0D#),
      3509 => to_slv(opcode_type, 16#0D#),
      3510 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#08#),
      3521 => to_slv(opcode_type, 16#05#),
      3522 => to_slv(opcode_type, 16#09#),
      3523 => to_slv(opcode_type, 16#06#),
      3524 => to_slv(opcode_type, 16#10#),
      3525 => to_slv(opcode_type, 16#0C#),
      3526 => to_slv(opcode_type, 16#05#),
      3527 => to_slv(opcode_type, 16#0A#),
      3528 => to_slv(opcode_type, 16#08#),
      3529 => to_slv(opcode_type, 16#08#),
      3530 => to_slv(opcode_type, 16#09#),
      3531 => to_slv(opcode_type, 16#10#),
      3532 => to_slv(opcode_type, 16#87#),
      3533 => to_slv(opcode_type, 16#08#),
      3534 => to_slv(opcode_type, 16#E2#),
      3535 => to_slv(opcode_type, 16#0A#),
      3536 => to_slv(opcode_type, 16#08#),
      3537 => to_slv(opcode_type, 16#09#),
      3538 => to_slv(opcode_type, 16#0A#),
      3539 => to_slv(opcode_type, 16#0E#),
      3540 => to_slv(opcode_type, 16#03#),
      3541 => to_slv(opcode_type, 16#0A#),
      3542 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#08#),
      3553 => to_slv(opcode_type, 16#08#),
      3554 => to_slv(opcode_type, 16#08#),
      3555 => to_slv(opcode_type, 16#07#),
      3556 => to_slv(opcode_type, 16#0A#),
      3557 => to_slv(opcode_type, 16#0F#),
      3558 => to_slv(opcode_type, 16#05#),
      3559 => to_slv(opcode_type, 16#0F#),
      3560 => to_slv(opcode_type, 16#08#),
      3561 => to_slv(opcode_type, 16#03#),
      3562 => to_slv(opcode_type, 16#0C#),
      3563 => to_slv(opcode_type, 16#03#),
      3564 => to_slv(opcode_type, 16#0C#),
      3565 => to_slv(opcode_type, 16#09#),
      3566 => to_slv(opcode_type, 16#02#),
      3567 => to_slv(opcode_type, 16#01#),
      3568 => to_slv(opcode_type, 16#0E#),
      3569 => to_slv(opcode_type, 16#08#),
      3570 => to_slv(opcode_type, 16#04#),
      3571 => to_slv(opcode_type, 16#0A#),
      3572 => to_slv(opcode_type, 16#02#),
      3573 => to_slv(opcode_type, 16#10#),
      3574 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#06#),
      3585 => to_slv(opcode_type, 16#02#),
      3586 => to_slv(opcode_type, 16#09#),
      3587 => to_slv(opcode_type, 16#08#),
      3588 => to_slv(opcode_type, 16#0D#),
      3589 => to_slv(opcode_type, 16#11#),
      3590 => to_slv(opcode_type, 16#06#),
      3591 => to_slv(opcode_type, 16#11#),
      3592 => to_slv(opcode_type, 16#0D#),
      3593 => to_slv(opcode_type, 16#06#),
      3594 => to_slv(opcode_type, 16#08#),
      3595 => to_slv(opcode_type, 16#09#),
      3596 => to_slv(opcode_type, 16#0C#),
      3597 => to_slv(opcode_type, 16#0C#),
      3598 => to_slv(opcode_type, 16#02#),
      3599 => to_slv(opcode_type, 16#0A#),
      3600 => to_slv(opcode_type, 16#08#),
      3601 => to_slv(opcode_type, 16#07#),
      3602 => to_slv(opcode_type, 16#0C#),
      3603 => to_slv(opcode_type, 16#0A#),
      3604 => to_slv(opcode_type, 16#02#),
      3605 => to_slv(opcode_type, 16#0C#),
      3606 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#07#),
      3617 => to_slv(opcode_type, 16#02#),
      3618 => to_slv(opcode_type, 16#07#),
      3619 => to_slv(opcode_type, 16#08#),
      3620 => to_slv(opcode_type, 16#5C#),
      3621 => to_slv(opcode_type, 16#11#),
      3622 => to_slv(opcode_type, 16#01#),
      3623 => to_slv(opcode_type, 16#0C#),
      3624 => to_slv(opcode_type, 16#09#),
      3625 => to_slv(opcode_type, 16#09#),
      3626 => to_slv(opcode_type, 16#07#),
      3627 => to_slv(opcode_type, 16#0E#),
      3628 => to_slv(opcode_type, 16#0B#),
      3629 => to_slv(opcode_type, 16#03#),
      3630 => to_slv(opcode_type, 16#0A#),
      3631 => to_slv(opcode_type, 16#07#),
      3632 => to_slv(opcode_type, 16#07#),
      3633 => to_slv(opcode_type, 16#0C#),
      3634 => to_slv(opcode_type, 16#0D#),
      3635 => to_slv(opcode_type, 16#09#),
      3636 => to_slv(opcode_type, 16#10#),
      3637 => to_slv(opcode_type, 16#0B#),
      3638 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#06#),
      3649 => to_slv(opcode_type, 16#09#),
      3650 => to_slv(opcode_type, 16#04#),
      3651 => to_slv(opcode_type, 16#04#),
      3652 => to_slv(opcode_type, 16#0E#),
      3653 => to_slv(opcode_type, 16#07#),
      3654 => to_slv(opcode_type, 16#01#),
      3655 => to_slv(opcode_type, 16#D9#),
      3656 => to_slv(opcode_type, 16#01#),
      3657 => to_slv(opcode_type, 16#10#),
      3658 => to_slv(opcode_type, 16#06#),
      3659 => to_slv(opcode_type, 16#08#),
      3660 => to_slv(opcode_type, 16#03#),
      3661 => to_slv(opcode_type, 16#0B#),
      3662 => to_slv(opcode_type, 16#04#),
      3663 => to_slv(opcode_type, 16#7B#),
      3664 => to_slv(opcode_type, 16#06#),
      3665 => to_slv(opcode_type, 16#03#),
      3666 => to_slv(opcode_type, 16#0B#),
      3667 => to_slv(opcode_type, 16#09#),
      3668 => to_slv(opcode_type, 16#0C#),
      3669 => to_slv(opcode_type, 16#10#),
      3670 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#06#),
      3681 => to_slv(opcode_type, 16#09#),
      3682 => to_slv(opcode_type, 16#05#),
      3683 => to_slv(opcode_type, 16#02#),
      3684 => to_slv(opcode_type, 16#0E#),
      3685 => to_slv(opcode_type, 16#04#),
      3686 => to_slv(opcode_type, 16#04#),
      3687 => to_slv(opcode_type, 16#0A#),
      3688 => to_slv(opcode_type, 16#08#),
      3689 => to_slv(opcode_type, 16#08#),
      3690 => to_slv(opcode_type, 16#05#),
      3691 => to_slv(opcode_type, 16#0B#),
      3692 => to_slv(opcode_type, 16#09#),
      3693 => to_slv(opcode_type, 16#0D#),
      3694 => to_slv(opcode_type, 16#0D#),
      3695 => to_slv(opcode_type, 16#06#),
      3696 => to_slv(opcode_type, 16#06#),
      3697 => to_slv(opcode_type, 16#0E#),
      3698 => to_slv(opcode_type, 16#0C#),
      3699 => to_slv(opcode_type, 16#07#),
      3700 => to_slv(opcode_type, 16#0B#),
      3701 => to_slv(opcode_type, 16#11#),
      3702 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#09#),
      3713 => to_slv(opcode_type, 16#02#),
      3714 => to_slv(opcode_type, 16#07#),
      3715 => to_slv(opcode_type, 16#03#),
      3716 => to_slv(opcode_type, 16#0D#),
      3717 => to_slv(opcode_type, 16#05#),
      3718 => to_slv(opcode_type, 16#FD#),
      3719 => to_slv(opcode_type, 16#06#),
      3720 => to_slv(opcode_type, 16#07#),
      3721 => to_slv(opcode_type, 16#09#),
      3722 => to_slv(opcode_type, 16#0E#),
      3723 => to_slv(opcode_type, 16#0D#),
      3724 => to_slv(opcode_type, 16#08#),
      3725 => to_slv(opcode_type, 16#A2#),
      3726 => to_slv(opcode_type, 16#0A#),
      3727 => to_slv(opcode_type, 16#08#),
      3728 => to_slv(opcode_type, 16#06#),
      3729 => to_slv(opcode_type, 16#11#),
      3730 => to_slv(opcode_type, 16#0A#),
      3731 => to_slv(opcode_type, 16#09#),
      3732 => to_slv(opcode_type, 16#C8#),
      3733 => to_slv(opcode_type, 16#42#),
      3734 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#07#),
      3745 => to_slv(opcode_type, 16#01#),
      3746 => to_slv(opcode_type, 16#07#),
      3747 => to_slv(opcode_type, 16#03#),
      3748 => to_slv(opcode_type, 16#0F#),
      3749 => to_slv(opcode_type, 16#05#),
      3750 => to_slv(opcode_type, 16#0E#),
      3751 => to_slv(opcode_type, 16#07#),
      3752 => to_slv(opcode_type, 16#09#),
      3753 => to_slv(opcode_type, 16#09#),
      3754 => to_slv(opcode_type, 16#5E#),
      3755 => to_slv(opcode_type, 16#0F#),
      3756 => to_slv(opcode_type, 16#06#),
      3757 => to_slv(opcode_type, 16#0C#),
      3758 => to_slv(opcode_type, 16#0A#),
      3759 => to_slv(opcode_type, 16#09#),
      3760 => to_slv(opcode_type, 16#07#),
      3761 => to_slv(opcode_type, 16#10#),
      3762 => to_slv(opcode_type, 16#0F#),
      3763 => to_slv(opcode_type, 16#07#),
      3764 => to_slv(opcode_type, 16#0C#),
      3765 => to_slv(opcode_type, 16#0E#),
      3766 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#08#),
      3777 => to_slv(opcode_type, 16#04#),
      3778 => to_slv(opcode_type, 16#09#),
      3779 => to_slv(opcode_type, 16#02#),
      3780 => to_slv(opcode_type, 16#11#),
      3781 => to_slv(opcode_type, 16#03#),
      3782 => to_slv(opcode_type, 16#0B#),
      3783 => to_slv(opcode_type, 16#06#),
      3784 => to_slv(opcode_type, 16#09#),
      3785 => to_slv(opcode_type, 16#06#),
      3786 => to_slv(opcode_type, 16#0C#),
      3787 => to_slv(opcode_type, 16#0A#),
      3788 => to_slv(opcode_type, 16#06#),
      3789 => to_slv(opcode_type, 16#0A#),
      3790 => to_slv(opcode_type, 16#10#),
      3791 => to_slv(opcode_type, 16#07#),
      3792 => to_slv(opcode_type, 16#07#),
      3793 => to_slv(opcode_type, 16#0C#),
      3794 => to_slv(opcode_type, 16#0D#),
      3795 => to_slv(opcode_type, 16#06#),
      3796 => to_slv(opcode_type, 16#0E#),
      3797 => to_slv(opcode_type, 16#0E#),
      3798 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#07#),
      3809 => to_slv(opcode_type, 16#04#),
      3810 => to_slv(opcode_type, 16#07#),
      3811 => to_slv(opcode_type, 16#06#),
      3812 => to_slv(opcode_type, 16#0D#),
      3813 => to_slv(opcode_type, 16#0F#),
      3814 => to_slv(opcode_type, 16#04#),
      3815 => to_slv(opcode_type, 16#0A#),
      3816 => to_slv(opcode_type, 16#09#),
      3817 => to_slv(opcode_type, 16#08#),
      3818 => to_slv(opcode_type, 16#03#),
      3819 => to_slv(opcode_type, 16#11#),
      3820 => to_slv(opcode_type, 16#09#),
      3821 => to_slv(opcode_type, 16#0B#),
      3822 => to_slv(opcode_type, 16#0F#),
      3823 => to_slv(opcode_type, 16#07#),
      3824 => to_slv(opcode_type, 16#09#),
      3825 => to_slv(opcode_type, 16#0B#),
      3826 => to_slv(opcode_type, 16#96#),
      3827 => to_slv(opcode_type, 16#09#),
      3828 => to_slv(opcode_type, 16#0B#),
      3829 => to_slv(opcode_type, 16#E6#),
      3830 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#06#),
      3841 => to_slv(opcode_type, 16#01#),
      3842 => to_slv(opcode_type, 16#07#),
      3843 => to_slv(opcode_type, 16#09#),
      3844 => to_slv(opcode_type, 16#0C#),
      3845 => to_slv(opcode_type, 16#0A#),
      3846 => to_slv(opcode_type, 16#02#),
      3847 => to_slv(opcode_type, 16#1D#),
      3848 => to_slv(opcode_type, 16#08#),
      3849 => to_slv(opcode_type, 16#06#),
      3850 => to_slv(opcode_type, 16#09#),
      3851 => to_slv(opcode_type, 16#0F#),
      3852 => to_slv(opcode_type, 16#9C#),
      3853 => to_slv(opcode_type, 16#01#),
      3854 => to_slv(opcode_type, 16#10#),
      3855 => to_slv(opcode_type, 16#06#),
      3856 => to_slv(opcode_type, 16#09#),
      3857 => to_slv(opcode_type, 16#10#),
      3858 => to_slv(opcode_type, 16#0D#),
      3859 => to_slv(opcode_type, 16#09#),
      3860 => to_slv(opcode_type, 16#0B#),
      3861 => to_slv(opcode_type, 16#38#),
      3862 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#07#),
      3873 => to_slv(opcode_type, 16#07#),
      3874 => to_slv(opcode_type, 16#03#),
      3875 => to_slv(opcode_type, 16#08#),
      3876 => to_slv(opcode_type, 16#11#),
      3877 => to_slv(opcode_type, 16#17#),
      3878 => to_slv(opcode_type, 16#09#),
      3879 => to_slv(opcode_type, 16#03#),
      3880 => to_slv(opcode_type, 16#10#),
      3881 => to_slv(opcode_type, 16#09#),
      3882 => to_slv(opcode_type, 16#0B#),
      3883 => to_slv(opcode_type, 16#0B#),
      3884 => to_slv(opcode_type, 16#06#),
      3885 => to_slv(opcode_type, 16#01#),
      3886 => to_slv(opcode_type, 16#01#),
      3887 => to_slv(opcode_type, 16#0A#),
      3888 => to_slv(opcode_type, 16#09#),
      3889 => to_slv(opcode_type, 16#01#),
      3890 => to_slv(opcode_type, 16#10#),
      3891 => to_slv(opcode_type, 16#07#),
      3892 => to_slv(opcode_type, 16#0D#),
      3893 => to_slv(opcode_type, 16#10#),
      3894 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#07#),
      3905 => to_slv(opcode_type, 16#05#),
      3906 => to_slv(opcode_type, 16#07#),
      3907 => to_slv(opcode_type, 16#04#),
      3908 => to_slv(opcode_type, 16#11#),
      3909 => to_slv(opcode_type, 16#09#),
      3910 => to_slv(opcode_type, 16#0A#),
      3911 => to_slv(opcode_type, 16#11#),
      3912 => to_slv(opcode_type, 16#07#),
      3913 => to_slv(opcode_type, 16#07#),
      3914 => to_slv(opcode_type, 16#07#),
      3915 => to_slv(opcode_type, 16#0A#),
      3916 => to_slv(opcode_type, 16#F9#),
      3917 => to_slv(opcode_type, 16#09#),
      3918 => to_slv(opcode_type, 16#0D#),
      3919 => to_slv(opcode_type, 16#8E#),
      3920 => to_slv(opcode_type, 16#09#),
      3921 => to_slv(opcode_type, 16#09#),
      3922 => to_slv(opcode_type, 16#10#),
      3923 => to_slv(opcode_type, 16#10#),
      3924 => to_slv(opcode_type, 16#03#),
      3925 => to_slv(opcode_type, 16#0F#),
      3926 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#07#),
      3937 => to_slv(opcode_type, 16#06#),
      3938 => to_slv(opcode_type, 16#07#),
      3939 => to_slv(opcode_type, 16#08#),
      3940 => to_slv(opcode_type, 16#0E#),
      3941 => to_slv(opcode_type, 16#11#),
      3942 => to_slv(opcode_type, 16#07#),
      3943 => to_slv(opcode_type, 16#0B#),
      3944 => to_slv(opcode_type, 16#26#),
      3945 => to_slv(opcode_type, 16#03#),
      3946 => to_slv(opcode_type, 16#07#),
      3947 => to_slv(opcode_type, 16#10#),
      3948 => to_slv(opcode_type, 16#0F#),
      3949 => to_slv(opcode_type, 16#06#),
      3950 => to_slv(opcode_type, 16#02#),
      3951 => to_slv(opcode_type, 16#05#),
      3952 => to_slv(opcode_type, 16#10#),
      3953 => to_slv(opcode_type, 16#06#),
      3954 => to_slv(opcode_type, 16#01#),
      3955 => to_slv(opcode_type, 16#0B#),
      3956 => to_slv(opcode_type, 16#05#),
      3957 => to_slv(opcode_type, 16#0D#),
      3958 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#06#),
      3969 => to_slv(opcode_type, 16#05#),
      3970 => to_slv(opcode_type, 16#09#),
      3971 => to_slv(opcode_type, 16#09#),
      3972 => to_slv(opcode_type, 16#11#),
      3973 => to_slv(opcode_type, 16#0A#),
      3974 => to_slv(opcode_type, 16#08#),
      3975 => to_slv(opcode_type, 16#0E#),
      3976 => to_slv(opcode_type, 16#0F#),
      3977 => to_slv(opcode_type, 16#09#),
      3978 => to_slv(opcode_type, 16#08#),
      3979 => to_slv(opcode_type, 16#04#),
      3980 => to_slv(opcode_type, 16#0A#),
      3981 => to_slv(opcode_type, 16#05#),
      3982 => to_slv(opcode_type, 16#0D#),
      3983 => to_slv(opcode_type, 16#09#),
      3984 => to_slv(opcode_type, 16#09#),
      3985 => to_slv(opcode_type, 16#FC#),
      3986 => to_slv(opcode_type, 16#0E#),
      3987 => to_slv(opcode_type, 16#06#),
      3988 => to_slv(opcode_type, 16#10#),
      3989 => to_slv(opcode_type, 16#10#),
      3990 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#06#),
      4001 => to_slv(opcode_type, 16#07#),
      4002 => to_slv(opcode_type, 16#08#),
      4003 => to_slv(opcode_type, 16#09#),
      4004 => to_slv(opcode_type, 16#0B#),
      4005 => to_slv(opcode_type, 16#0F#),
      4006 => to_slv(opcode_type, 16#05#),
      4007 => to_slv(opcode_type, 16#0F#),
      4008 => to_slv(opcode_type, 16#02#),
      4009 => to_slv(opcode_type, 16#06#),
      4010 => to_slv(opcode_type, 16#11#),
      4011 => to_slv(opcode_type, 16#0F#),
      4012 => to_slv(opcode_type, 16#08#),
      4013 => to_slv(opcode_type, 16#07#),
      4014 => to_slv(opcode_type, 16#07#),
      4015 => to_slv(opcode_type, 16#0C#),
      4016 => to_slv(opcode_type, 16#0E#),
      4017 => to_slv(opcode_type, 16#05#),
      4018 => to_slv(opcode_type, 16#0B#),
      4019 => to_slv(opcode_type, 16#02#),
      4020 => to_slv(opcode_type, 16#05#),
      4021 => to_slv(opcode_type, 16#8A#),
      4022 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#07#),
      4033 => to_slv(opcode_type, 16#04#),
      4034 => to_slv(opcode_type, 16#08#),
      4035 => to_slv(opcode_type, 16#08#),
      4036 => to_slv(opcode_type, 16#0F#),
      4037 => to_slv(opcode_type, 16#10#),
      4038 => to_slv(opcode_type, 16#04#),
      4039 => to_slv(opcode_type, 16#10#),
      4040 => to_slv(opcode_type, 16#09#),
      4041 => to_slv(opcode_type, 16#06#),
      4042 => to_slv(opcode_type, 16#01#),
      4043 => to_slv(opcode_type, 16#0F#),
      4044 => to_slv(opcode_type, 16#07#),
      4045 => to_slv(opcode_type, 16#0C#),
      4046 => to_slv(opcode_type, 16#82#),
      4047 => to_slv(opcode_type, 16#08#),
      4048 => to_slv(opcode_type, 16#06#),
      4049 => to_slv(opcode_type, 16#11#),
      4050 => to_slv(opcode_type, 16#0F#),
      4051 => to_slv(opcode_type, 16#06#),
      4052 => to_slv(opcode_type, 16#0E#),
      4053 => to_slv(opcode_type, 16#0D#),
      4054 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#08#),
      4065 => to_slv(opcode_type, 16#08#),
      4066 => to_slv(opcode_type, 16#04#),
      4067 => to_slv(opcode_type, 16#02#),
      4068 => to_slv(opcode_type, 16#0F#),
      4069 => to_slv(opcode_type, 16#04#),
      4070 => to_slv(opcode_type, 16#09#),
      4071 => to_slv(opcode_type, 16#10#),
      4072 => to_slv(opcode_type, 16#0B#),
      4073 => to_slv(opcode_type, 16#06#),
      4074 => to_slv(opcode_type, 16#09#),
      4075 => to_slv(opcode_type, 16#05#),
      4076 => to_slv(opcode_type, 16#0E#),
      4077 => to_slv(opcode_type, 16#09#),
      4078 => to_slv(opcode_type, 16#0B#),
      4079 => to_slv(opcode_type, 16#0E#),
      4080 => to_slv(opcode_type, 16#07#),
      4081 => to_slv(opcode_type, 16#07#),
      4082 => to_slv(opcode_type, 16#0C#),
      4083 => to_slv(opcode_type, 16#10#),
      4084 => to_slv(opcode_type, 16#04#),
      4085 => to_slv(opcode_type, 16#0E#),
      4086 to 4095 => (others => '0')
  ),

    -- Bin `23`...
    22 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#08#),
      1 => to_slv(opcode_type, 16#06#),
      2 => to_slv(opcode_type, 16#02#),
      3 => to_slv(opcode_type, 16#04#),
      4 => to_slv(opcode_type, 16#0B#),
      5 => to_slv(opcode_type, 16#04#),
      6 => to_slv(opcode_type, 16#07#),
      7 => to_slv(opcode_type, 16#10#),
      8 => to_slv(opcode_type, 16#0D#),
      9 => to_slv(opcode_type, 16#06#),
      10 => to_slv(opcode_type, 16#07#),
      11 => to_slv(opcode_type, 16#01#),
      12 => to_slv(opcode_type, 16#10#),
      13 => to_slv(opcode_type, 16#09#),
      14 => to_slv(opcode_type, 16#0A#),
      15 => to_slv(opcode_type, 16#0E#),
      16 => to_slv(opcode_type, 16#07#),
      17 => to_slv(opcode_type, 16#06#),
      18 => to_slv(opcode_type, 16#0B#),
      19 => to_slv(opcode_type, 16#11#),
      20 => to_slv(opcode_type, 16#09#),
      21 => to_slv(opcode_type, 16#0A#),
      22 => to_slv(opcode_type, 16#0B#),
      23 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#09#),
      33 => to_slv(opcode_type, 16#09#),
      34 => to_slv(opcode_type, 16#02#),
      35 => to_slv(opcode_type, 16#03#),
      36 => to_slv(opcode_type, 16#0E#),
      37 => to_slv(opcode_type, 16#03#),
      38 => to_slv(opcode_type, 16#01#),
      39 => to_slv(opcode_type, 16#FB#),
      40 => to_slv(opcode_type, 16#06#),
      41 => to_slv(opcode_type, 16#09#),
      42 => to_slv(opcode_type, 16#06#),
      43 => to_slv(opcode_type, 16#0C#),
      44 => to_slv(opcode_type, 16#0A#),
      45 => to_slv(opcode_type, 16#09#),
      46 => to_slv(opcode_type, 16#0A#),
      47 => to_slv(opcode_type, 16#37#),
      48 => to_slv(opcode_type, 16#06#),
      49 => to_slv(opcode_type, 16#07#),
      50 => to_slv(opcode_type, 16#0F#),
      51 => to_slv(opcode_type, 16#0F#),
      52 => to_slv(opcode_type, 16#06#),
      53 => to_slv(opcode_type, 16#0F#),
      54 => to_slv(opcode_type, 16#0B#),
      55 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#08#),
      65 => to_slv(opcode_type, 16#02#),
      66 => to_slv(opcode_type, 16#07#),
      67 => to_slv(opcode_type, 16#04#),
      68 => to_slv(opcode_type, 16#0B#),
      69 => to_slv(opcode_type, 16#08#),
      70 => to_slv(opcode_type, 16#11#),
      71 => to_slv(opcode_type, 16#0F#),
      72 => to_slv(opcode_type, 16#06#),
      73 => to_slv(opcode_type, 16#08#),
      74 => to_slv(opcode_type, 16#07#),
      75 => to_slv(opcode_type, 16#0A#),
      76 => to_slv(opcode_type, 16#0D#),
      77 => to_slv(opcode_type, 16#08#),
      78 => to_slv(opcode_type, 16#0E#),
      79 => to_slv(opcode_type, 16#0B#),
      80 => to_slv(opcode_type, 16#09#),
      81 => to_slv(opcode_type, 16#08#),
      82 => to_slv(opcode_type, 16#10#),
      83 => to_slv(opcode_type, 16#0A#),
      84 => to_slv(opcode_type, 16#06#),
      85 => to_slv(opcode_type, 16#0A#),
      86 => to_slv(opcode_type, 16#0E#),
      87 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#06#),
      97 => to_slv(opcode_type, 16#02#),
      98 => to_slv(opcode_type, 16#09#),
      99 => to_slv(opcode_type, 16#05#),
      100 => to_slv(opcode_type, 16#0A#),
      101 => to_slv(opcode_type, 16#08#),
      102 => to_slv(opcode_type, 16#0C#),
      103 => to_slv(opcode_type, 16#0B#),
      104 => to_slv(opcode_type, 16#07#),
      105 => to_slv(opcode_type, 16#07#),
      106 => to_slv(opcode_type, 16#08#),
      107 => to_slv(opcode_type, 16#0C#),
      108 => to_slv(opcode_type, 16#0D#),
      109 => to_slv(opcode_type, 16#09#),
      110 => to_slv(opcode_type, 16#0A#),
      111 => to_slv(opcode_type, 16#11#),
      112 => to_slv(opcode_type, 16#09#),
      113 => to_slv(opcode_type, 16#07#),
      114 => to_slv(opcode_type, 16#0C#),
      115 => to_slv(opcode_type, 16#10#),
      116 => to_slv(opcode_type, 16#06#),
      117 => to_slv(opcode_type, 16#0D#),
      118 => to_slv(opcode_type, 16#0F#),
      119 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#08#),
      129 => to_slv(opcode_type, 16#08#),
      130 => to_slv(opcode_type, 16#05#),
      131 => to_slv(opcode_type, 16#07#),
      132 => to_slv(opcode_type, 16#11#),
      133 => to_slv(opcode_type, 16#0C#),
      134 => to_slv(opcode_type, 16#08#),
      135 => to_slv(opcode_type, 16#05#),
      136 => to_slv(opcode_type, 16#0D#),
      137 => to_slv(opcode_type, 16#07#),
      138 => to_slv(opcode_type, 16#0E#),
      139 => to_slv(opcode_type, 16#0C#),
      140 => to_slv(opcode_type, 16#08#),
      141 => to_slv(opcode_type, 16#08#),
      142 => to_slv(opcode_type, 16#06#),
      143 => to_slv(opcode_type, 16#4C#),
      144 => to_slv(opcode_type, 16#0F#),
      145 => to_slv(opcode_type, 16#02#),
      146 => to_slv(opcode_type, 16#0C#),
      147 => to_slv(opcode_type, 16#01#),
      148 => to_slv(opcode_type, 16#07#),
      149 => to_slv(opcode_type, 16#0F#),
      150 => to_slv(opcode_type, 16#0C#),
      151 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#07#),
      161 => to_slv(opcode_type, 16#01#),
      162 => to_slv(opcode_type, 16#06#),
      163 => to_slv(opcode_type, 16#04#),
      164 => to_slv(opcode_type, 16#6B#),
      165 => to_slv(opcode_type, 16#09#),
      166 => to_slv(opcode_type, 16#0D#),
      167 => to_slv(opcode_type, 16#0B#),
      168 => to_slv(opcode_type, 16#09#),
      169 => to_slv(opcode_type, 16#09#),
      170 => to_slv(opcode_type, 16#07#),
      171 => to_slv(opcode_type, 16#0A#),
      172 => to_slv(opcode_type, 16#0D#),
      173 => to_slv(opcode_type, 16#08#),
      174 => to_slv(opcode_type, 16#10#),
      175 => to_slv(opcode_type, 16#11#),
      176 => to_slv(opcode_type, 16#06#),
      177 => to_slv(opcode_type, 16#06#),
      178 => to_slv(opcode_type, 16#0E#),
      179 => to_slv(opcode_type, 16#0A#),
      180 => to_slv(opcode_type, 16#07#),
      181 => to_slv(opcode_type, 16#0D#),
      182 => to_slv(opcode_type, 16#10#),
      183 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#09#),
      193 => to_slv(opcode_type, 16#08#),
      194 => to_slv(opcode_type, 16#05#),
      195 => to_slv(opcode_type, 16#03#),
      196 => to_slv(opcode_type, 16#0D#),
      197 => to_slv(opcode_type, 16#03#),
      198 => to_slv(opcode_type, 16#06#),
      199 => to_slv(opcode_type, 16#0B#),
      200 => to_slv(opcode_type, 16#0C#),
      201 => to_slv(opcode_type, 16#08#),
      202 => to_slv(opcode_type, 16#06#),
      203 => to_slv(opcode_type, 16#02#),
      204 => to_slv(opcode_type, 16#0C#),
      205 => to_slv(opcode_type, 16#06#),
      206 => to_slv(opcode_type, 16#C7#),
      207 => to_slv(opcode_type, 16#0F#),
      208 => to_slv(opcode_type, 16#07#),
      209 => to_slv(opcode_type, 16#08#),
      210 => to_slv(opcode_type, 16#0D#),
      211 => to_slv(opcode_type, 16#10#),
      212 => to_slv(opcode_type, 16#08#),
      213 => to_slv(opcode_type, 16#0E#),
      214 => to_slv(opcode_type, 16#0A#),
      215 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#06#),
      225 => to_slv(opcode_type, 16#06#),
      226 => to_slv(opcode_type, 16#01#),
      227 => to_slv(opcode_type, 16#06#),
      228 => to_slv(opcode_type, 16#0C#),
      229 => to_slv(opcode_type, 16#10#),
      230 => to_slv(opcode_type, 16#09#),
      231 => to_slv(opcode_type, 16#05#),
      232 => to_slv(opcode_type, 16#10#),
      233 => to_slv(opcode_type, 16#05#),
      234 => to_slv(opcode_type, 16#0B#),
      235 => to_slv(opcode_type, 16#09#),
      236 => to_slv(opcode_type, 16#04#),
      237 => to_slv(opcode_type, 16#07#),
      238 => to_slv(opcode_type, 16#0B#),
      239 => to_slv(opcode_type, 16#0A#),
      240 => to_slv(opcode_type, 16#08#),
      241 => to_slv(opcode_type, 16#06#),
      242 => to_slv(opcode_type, 16#0D#),
      243 => to_slv(opcode_type, 16#0F#),
      244 => to_slv(opcode_type, 16#07#),
      245 => to_slv(opcode_type, 16#10#),
      246 => to_slv(opcode_type, 16#0A#),
      247 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#06#),
      257 => to_slv(opcode_type, 16#08#),
      258 => to_slv(opcode_type, 16#04#),
      259 => to_slv(opcode_type, 16#05#),
      260 => to_slv(opcode_type, 16#0F#),
      261 => to_slv(opcode_type, 16#08#),
      262 => to_slv(opcode_type, 16#09#),
      263 => to_slv(opcode_type, 16#0E#),
      264 => to_slv(opcode_type, 16#10#),
      265 => to_slv(opcode_type, 16#07#),
      266 => to_slv(opcode_type, 16#0A#),
      267 => to_slv(opcode_type, 16#10#),
      268 => to_slv(opcode_type, 16#09#),
      269 => to_slv(opcode_type, 16#03#),
      270 => to_slv(opcode_type, 16#02#),
      271 => to_slv(opcode_type, 16#10#),
      272 => to_slv(opcode_type, 16#08#),
      273 => to_slv(opcode_type, 16#06#),
      274 => to_slv(opcode_type, 16#0C#),
      275 => to_slv(opcode_type, 16#0D#),
      276 => to_slv(opcode_type, 16#08#),
      277 => to_slv(opcode_type, 16#5C#),
      278 => to_slv(opcode_type, 16#0B#),
      279 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#07#),
      290 => to_slv(opcode_type, 16#09#),
      291 => to_slv(opcode_type, 16#03#),
      292 => to_slv(opcode_type, 16#11#),
      293 => to_slv(opcode_type, 16#01#),
      294 => to_slv(opcode_type, 16#0A#),
      295 => to_slv(opcode_type, 16#06#),
      296 => to_slv(opcode_type, 16#01#),
      297 => to_slv(opcode_type, 16#0D#),
      298 => to_slv(opcode_type, 16#03#),
      299 => to_slv(opcode_type, 16#0E#),
      300 => to_slv(opcode_type, 16#08#),
      301 => to_slv(opcode_type, 16#06#),
      302 => to_slv(opcode_type, 16#04#),
      303 => to_slv(opcode_type, 16#0C#),
      304 => to_slv(opcode_type, 16#02#),
      305 => to_slv(opcode_type, 16#0A#),
      306 => to_slv(opcode_type, 16#06#),
      307 => to_slv(opcode_type, 16#09#),
      308 => to_slv(opcode_type, 16#0C#),
      309 => to_slv(opcode_type, 16#0B#),
      310 => to_slv(opcode_type, 16#B6#),
      311 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#06#),
      321 => to_slv(opcode_type, 16#01#),
      322 => to_slv(opcode_type, 16#09#),
      323 => to_slv(opcode_type, 16#05#),
      324 => to_slv(opcode_type, 16#0C#),
      325 => to_slv(opcode_type, 16#08#),
      326 => to_slv(opcode_type, 16#0A#),
      327 => to_slv(opcode_type, 16#0E#),
      328 => to_slv(opcode_type, 16#07#),
      329 => to_slv(opcode_type, 16#09#),
      330 => to_slv(opcode_type, 16#09#),
      331 => to_slv(opcode_type, 16#67#),
      332 => to_slv(opcode_type, 16#E5#),
      333 => to_slv(opcode_type, 16#06#),
      334 => to_slv(opcode_type, 16#0A#),
      335 => to_slv(opcode_type, 16#0A#),
      336 => to_slv(opcode_type, 16#06#),
      337 => to_slv(opcode_type, 16#06#),
      338 => to_slv(opcode_type, 16#0A#),
      339 => to_slv(opcode_type, 16#CA#),
      340 => to_slv(opcode_type, 16#08#),
      341 => to_slv(opcode_type, 16#10#),
      342 => to_slv(opcode_type, 16#11#),
      343 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#07#),
      353 => to_slv(opcode_type, 16#03#),
      354 => to_slv(opcode_type, 16#09#),
      355 => to_slv(opcode_type, 16#08#),
      356 => to_slv(opcode_type, 16#11#),
      357 => to_slv(opcode_type, 16#0C#),
      358 => to_slv(opcode_type, 16#03#),
      359 => to_slv(opcode_type, 16#1C#),
      360 => to_slv(opcode_type, 16#06#),
      361 => to_slv(opcode_type, 16#06#),
      362 => to_slv(opcode_type, 16#08#),
      363 => to_slv(opcode_type, 16#0A#),
      364 => to_slv(opcode_type, 16#0D#),
      365 => to_slv(opcode_type, 16#08#),
      366 => to_slv(opcode_type, 16#0A#),
      367 => to_slv(opcode_type, 16#AF#),
      368 => to_slv(opcode_type, 16#06#),
      369 => to_slv(opcode_type, 16#08#),
      370 => to_slv(opcode_type, 16#0D#),
      371 => to_slv(opcode_type, 16#0C#),
      372 => to_slv(opcode_type, 16#06#),
      373 => to_slv(opcode_type, 16#0E#),
      374 => to_slv(opcode_type, 16#11#),
      375 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#09#),
      385 => to_slv(opcode_type, 16#01#),
      386 => to_slv(opcode_type, 16#07#),
      387 => to_slv(opcode_type, 16#06#),
      388 => to_slv(opcode_type, 16#0B#),
      389 => to_slv(opcode_type, 16#0A#),
      390 => to_slv(opcode_type, 16#03#),
      391 => to_slv(opcode_type, 16#0F#),
      392 => to_slv(opcode_type, 16#09#),
      393 => to_slv(opcode_type, 16#07#),
      394 => to_slv(opcode_type, 16#07#),
      395 => to_slv(opcode_type, 16#0A#),
      396 => to_slv(opcode_type, 16#11#),
      397 => to_slv(opcode_type, 16#09#),
      398 => to_slv(opcode_type, 16#0A#),
      399 => to_slv(opcode_type, 16#10#),
      400 => to_slv(opcode_type, 16#08#),
      401 => to_slv(opcode_type, 16#08#),
      402 => to_slv(opcode_type, 16#0F#),
      403 => to_slv(opcode_type, 16#0A#),
      404 => to_slv(opcode_type, 16#09#),
      405 => to_slv(opcode_type, 16#0F#),
      406 => to_slv(opcode_type, 16#0D#),
      407 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#07#),
      417 => to_slv(opcode_type, 16#05#),
      418 => to_slv(opcode_type, 16#07#),
      419 => to_slv(opcode_type, 16#05#),
      420 => to_slv(opcode_type, 16#0F#),
      421 => to_slv(opcode_type, 16#06#),
      422 => to_slv(opcode_type, 16#10#),
      423 => to_slv(opcode_type, 16#0F#),
      424 => to_slv(opcode_type, 16#07#),
      425 => to_slv(opcode_type, 16#09#),
      426 => to_slv(opcode_type, 16#09#),
      427 => to_slv(opcode_type, 16#0D#),
      428 => to_slv(opcode_type, 16#0A#),
      429 => to_slv(opcode_type, 16#06#),
      430 => to_slv(opcode_type, 16#0C#),
      431 => to_slv(opcode_type, 16#D9#),
      432 => to_slv(opcode_type, 16#07#),
      433 => to_slv(opcode_type, 16#06#),
      434 => to_slv(opcode_type, 16#0E#),
      435 => to_slv(opcode_type, 16#10#),
      436 => to_slv(opcode_type, 16#07#),
      437 => to_slv(opcode_type, 16#0F#),
      438 => to_slv(opcode_type, 16#0C#),
      439 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#06#),
      449 => to_slv(opcode_type, 16#07#),
      450 => to_slv(opcode_type, 16#04#),
      451 => to_slv(opcode_type, 16#06#),
      452 => to_slv(opcode_type, 16#0B#),
      453 => to_slv(opcode_type, 16#0D#),
      454 => to_slv(opcode_type, 16#04#),
      455 => to_slv(opcode_type, 16#09#),
      456 => to_slv(opcode_type, 16#0D#),
      457 => to_slv(opcode_type, 16#6F#),
      458 => to_slv(opcode_type, 16#09#),
      459 => to_slv(opcode_type, 16#07#),
      460 => to_slv(opcode_type, 16#01#),
      461 => to_slv(opcode_type, 16#0F#),
      462 => to_slv(opcode_type, 16#04#),
      463 => to_slv(opcode_type, 16#0B#),
      464 => to_slv(opcode_type, 16#06#),
      465 => to_slv(opcode_type, 16#08#),
      466 => to_slv(opcode_type, 16#0E#),
      467 => to_slv(opcode_type, 16#0B#),
      468 => to_slv(opcode_type, 16#07#),
      469 => to_slv(opcode_type, 16#0C#),
      470 => to_slv(opcode_type, 16#0D#),
      471 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#09#),
      481 => to_slv(opcode_type, 16#05#),
      482 => to_slv(opcode_type, 16#08#),
      483 => to_slv(opcode_type, 16#02#),
      484 => to_slv(opcode_type, 16#0C#),
      485 => to_slv(opcode_type, 16#08#),
      486 => to_slv(opcode_type, 16#0D#),
      487 => to_slv(opcode_type, 16#11#),
      488 => to_slv(opcode_type, 16#09#),
      489 => to_slv(opcode_type, 16#07#),
      490 => to_slv(opcode_type, 16#09#),
      491 => to_slv(opcode_type, 16#0A#),
      492 => to_slv(opcode_type, 16#10#),
      493 => to_slv(opcode_type, 16#07#),
      494 => to_slv(opcode_type, 16#10#),
      495 => to_slv(opcode_type, 16#10#),
      496 => to_slv(opcode_type, 16#09#),
      497 => to_slv(opcode_type, 16#06#),
      498 => to_slv(opcode_type, 16#11#),
      499 => to_slv(opcode_type, 16#11#),
      500 => to_slv(opcode_type, 16#07#),
      501 => to_slv(opcode_type, 16#0A#),
      502 => to_slv(opcode_type, 16#10#),
      503 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#07#),
      513 => to_slv(opcode_type, 16#04#),
      514 => to_slv(opcode_type, 16#06#),
      515 => to_slv(opcode_type, 16#04#),
      516 => to_slv(opcode_type, 16#0F#),
      517 => to_slv(opcode_type, 16#07#),
      518 => to_slv(opcode_type, 16#0C#),
      519 => to_slv(opcode_type, 16#0E#),
      520 => to_slv(opcode_type, 16#07#),
      521 => to_slv(opcode_type, 16#08#),
      522 => to_slv(opcode_type, 16#09#),
      523 => to_slv(opcode_type, 16#0D#),
      524 => to_slv(opcode_type, 16#0E#),
      525 => to_slv(opcode_type, 16#07#),
      526 => to_slv(opcode_type, 16#0E#),
      527 => to_slv(opcode_type, 16#0C#),
      528 => to_slv(opcode_type, 16#09#),
      529 => to_slv(opcode_type, 16#06#),
      530 => to_slv(opcode_type, 16#0B#),
      531 => to_slv(opcode_type, 16#B6#),
      532 => to_slv(opcode_type, 16#06#),
      533 => to_slv(opcode_type, 16#0C#),
      534 => to_slv(opcode_type, 16#11#),
      535 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#07#),
      545 => to_slv(opcode_type, 16#06#),
      546 => to_slv(opcode_type, 16#06#),
      547 => to_slv(opcode_type, 16#06#),
      548 => to_slv(opcode_type, 16#B9#),
      549 => to_slv(opcode_type, 16#0E#),
      550 => to_slv(opcode_type, 16#09#),
      551 => to_slv(opcode_type, 16#0B#),
      552 => to_slv(opcode_type, 16#0C#),
      553 => to_slv(opcode_type, 16#01#),
      554 => to_slv(opcode_type, 16#03#),
      555 => to_slv(opcode_type, 16#0C#),
      556 => to_slv(opcode_type, 16#07#),
      557 => to_slv(opcode_type, 16#07#),
      558 => to_slv(opcode_type, 16#07#),
      559 => to_slv(opcode_type, 16#0D#),
      560 => to_slv(opcode_type, 16#0F#),
      561 => to_slv(opcode_type, 16#02#),
      562 => to_slv(opcode_type, 16#0E#),
      563 => to_slv(opcode_type, 16#07#),
      564 => to_slv(opcode_type, 16#04#),
      565 => to_slv(opcode_type, 16#10#),
      566 => to_slv(opcode_type, 16#0A#),
      567 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#09#),
      577 => to_slv(opcode_type, 16#01#),
      578 => to_slv(opcode_type, 16#09#),
      579 => to_slv(opcode_type, 16#04#),
      580 => to_slv(opcode_type, 16#0F#),
      581 => to_slv(opcode_type, 16#06#),
      582 => to_slv(opcode_type, 16#11#),
      583 => to_slv(opcode_type, 16#0E#),
      584 => to_slv(opcode_type, 16#08#),
      585 => to_slv(opcode_type, 16#09#),
      586 => to_slv(opcode_type, 16#09#),
      587 => to_slv(opcode_type, 16#0C#),
      588 => to_slv(opcode_type, 16#0A#),
      589 => to_slv(opcode_type, 16#06#),
      590 => to_slv(opcode_type, 16#0C#),
      591 => to_slv(opcode_type, 16#0C#),
      592 => to_slv(opcode_type, 16#06#),
      593 => to_slv(opcode_type, 16#09#),
      594 => to_slv(opcode_type, 16#0E#),
      595 => to_slv(opcode_type, 16#6E#),
      596 => to_slv(opcode_type, 16#07#),
      597 => to_slv(opcode_type, 16#0A#),
      598 => to_slv(opcode_type, 16#0F#),
      599 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#07#),
      609 => to_slv(opcode_type, 16#03#),
      610 => to_slv(opcode_type, 16#08#),
      611 => to_slv(opcode_type, 16#07#),
      612 => to_slv(opcode_type, 16#0E#),
      613 => to_slv(opcode_type, 16#11#),
      614 => to_slv(opcode_type, 16#01#),
      615 => to_slv(opcode_type, 16#EC#),
      616 => to_slv(opcode_type, 16#08#),
      617 => to_slv(opcode_type, 16#08#),
      618 => to_slv(opcode_type, 16#09#),
      619 => to_slv(opcode_type, 16#0D#),
      620 => to_slv(opcode_type, 16#0A#),
      621 => to_slv(opcode_type, 16#08#),
      622 => to_slv(opcode_type, 16#0F#),
      623 => to_slv(opcode_type, 16#0E#),
      624 => to_slv(opcode_type, 16#06#),
      625 => to_slv(opcode_type, 16#09#),
      626 => to_slv(opcode_type, 16#0B#),
      627 => to_slv(opcode_type, 16#0B#),
      628 => to_slv(opcode_type, 16#08#),
      629 => to_slv(opcode_type, 16#11#),
      630 => to_slv(opcode_type, 16#0E#),
      631 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#07#),
      641 => to_slv(opcode_type, 16#09#),
      642 => to_slv(opcode_type, 16#07#),
      643 => to_slv(opcode_type, 16#09#),
      644 => to_slv(opcode_type, 16#0E#),
      645 => to_slv(opcode_type, 16#0E#),
      646 => to_slv(opcode_type, 16#05#),
      647 => to_slv(opcode_type, 16#0E#),
      648 => to_slv(opcode_type, 16#03#),
      649 => to_slv(opcode_type, 16#08#),
      650 => to_slv(opcode_type, 16#0C#),
      651 => to_slv(opcode_type, 16#0A#),
      652 => to_slv(opcode_type, 16#08#),
      653 => to_slv(opcode_type, 16#09#),
      654 => to_slv(opcode_type, 16#07#),
      655 => to_slv(opcode_type, 16#0C#),
      656 => to_slv(opcode_type, 16#11#),
      657 => to_slv(opcode_type, 16#07#),
      658 => to_slv(opcode_type, 16#0E#),
      659 => to_slv(opcode_type, 16#0A#),
      660 => to_slv(opcode_type, 16#01#),
      661 => to_slv(opcode_type, 16#01#),
      662 => to_slv(opcode_type, 16#0A#),
      663 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#09#),
      673 => to_slv(opcode_type, 16#07#),
      674 => to_slv(opcode_type, 16#05#),
      675 => to_slv(opcode_type, 16#03#),
      676 => to_slv(opcode_type, 16#0B#),
      677 => to_slv(opcode_type, 16#08#),
      678 => to_slv(opcode_type, 16#03#),
      679 => to_slv(opcode_type, 16#0E#),
      680 => to_slv(opcode_type, 16#02#),
      681 => to_slv(opcode_type, 16#0E#),
      682 => to_slv(opcode_type, 16#09#),
      683 => to_slv(opcode_type, 16#07#),
      684 => to_slv(opcode_type, 16#02#),
      685 => to_slv(opcode_type, 16#A8#),
      686 => to_slv(opcode_type, 16#03#),
      687 => to_slv(opcode_type, 16#0F#),
      688 => to_slv(opcode_type, 16#08#),
      689 => to_slv(opcode_type, 16#08#),
      690 => to_slv(opcode_type, 16#0A#),
      691 => to_slv(opcode_type, 16#0C#),
      692 => to_slv(opcode_type, 16#09#),
      693 => to_slv(opcode_type, 16#10#),
      694 => to_slv(opcode_type, 16#0C#),
      695 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#08#),
      705 => to_slv(opcode_type, 16#03#),
      706 => to_slv(opcode_type, 16#06#),
      707 => to_slv(opcode_type, 16#02#),
      708 => to_slv(opcode_type, 16#0D#),
      709 => to_slv(opcode_type, 16#08#),
      710 => to_slv(opcode_type, 16#0B#),
      711 => to_slv(opcode_type, 16#11#),
      712 => to_slv(opcode_type, 16#09#),
      713 => to_slv(opcode_type, 16#09#),
      714 => to_slv(opcode_type, 16#07#),
      715 => to_slv(opcode_type, 16#0E#),
      716 => to_slv(opcode_type, 16#0E#),
      717 => to_slv(opcode_type, 16#06#),
      718 => to_slv(opcode_type, 16#0D#),
      719 => to_slv(opcode_type, 16#11#),
      720 => to_slv(opcode_type, 16#08#),
      721 => to_slv(opcode_type, 16#07#),
      722 => to_slv(opcode_type, 16#0F#),
      723 => to_slv(opcode_type, 16#0B#),
      724 => to_slv(opcode_type, 16#06#),
      725 => to_slv(opcode_type, 16#0D#),
      726 => to_slv(opcode_type, 16#0D#),
      727 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#08#),
      737 => to_slv(opcode_type, 16#04#),
      738 => to_slv(opcode_type, 16#07#),
      739 => to_slv(opcode_type, 16#06#),
      740 => to_slv(opcode_type, 16#0A#),
      741 => to_slv(opcode_type, 16#0F#),
      742 => to_slv(opcode_type, 16#04#),
      743 => to_slv(opcode_type, 16#11#),
      744 => to_slv(opcode_type, 16#08#),
      745 => to_slv(opcode_type, 16#08#),
      746 => to_slv(opcode_type, 16#08#),
      747 => to_slv(opcode_type, 16#10#),
      748 => to_slv(opcode_type, 16#0D#),
      749 => to_slv(opcode_type, 16#09#),
      750 => to_slv(opcode_type, 16#0D#),
      751 => to_slv(opcode_type, 16#0B#),
      752 => to_slv(opcode_type, 16#09#),
      753 => to_slv(opcode_type, 16#06#),
      754 => to_slv(opcode_type, 16#0A#),
      755 => to_slv(opcode_type, 16#10#),
      756 => to_slv(opcode_type, 16#06#),
      757 => to_slv(opcode_type, 16#11#),
      758 => to_slv(opcode_type, 16#0A#),
      759 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#06#),
      769 => to_slv(opcode_type, 16#08#),
      770 => to_slv(opcode_type, 16#04#),
      771 => to_slv(opcode_type, 16#01#),
      772 => to_slv(opcode_type, 16#0E#),
      773 => to_slv(opcode_type, 16#06#),
      774 => to_slv(opcode_type, 16#01#),
      775 => to_slv(opcode_type, 16#10#),
      776 => to_slv(opcode_type, 16#06#),
      777 => to_slv(opcode_type, 16#0F#),
      778 => to_slv(opcode_type, 16#0D#),
      779 => to_slv(opcode_type, 16#09#),
      780 => to_slv(opcode_type, 16#05#),
      781 => to_slv(opcode_type, 16#06#),
      782 => to_slv(opcode_type, 16#0B#),
      783 => to_slv(opcode_type, 16#0B#),
      784 => to_slv(opcode_type, 16#09#),
      785 => to_slv(opcode_type, 16#08#),
      786 => to_slv(opcode_type, 16#D3#),
      787 => to_slv(opcode_type, 16#0E#),
      788 => to_slv(opcode_type, 16#08#),
      789 => to_slv(opcode_type, 16#0A#),
      790 => to_slv(opcode_type, 16#0F#),
      791 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#06#),
      801 => to_slv(opcode_type, 16#04#),
      802 => to_slv(opcode_type, 16#09#),
      803 => to_slv(opcode_type, 16#02#),
      804 => to_slv(opcode_type, 16#0E#),
      805 => to_slv(opcode_type, 16#07#),
      806 => to_slv(opcode_type, 16#0E#),
      807 => to_slv(opcode_type, 16#0B#),
      808 => to_slv(opcode_type, 16#06#),
      809 => to_slv(opcode_type, 16#09#),
      810 => to_slv(opcode_type, 16#08#),
      811 => to_slv(opcode_type, 16#10#),
      812 => to_slv(opcode_type, 16#11#),
      813 => to_slv(opcode_type, 16#09#),
      814 => to_slv(opcode_type, 16#0C#),
      815 => to_slv(opcode_type, 16#D1#),
      816 => to_slv(opcode_type, 16#07#),
      817 => to_slv(opcode_type, 16#06#),
      818 => to_slv(opcode_type, 16#FF#),
      819 => to_slv(opcode_type, 16#0D#),
      820 => to_slv(opcode_type, 16#07#),
      821 => to_slv(opcode_type, 16#0F#),
      822 => to_slv(opcode_type, 16#0A#),
      823 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#08#),
      833 => to_slv(opcode_type, 16#01#),
      834 => to_slv(opcode_type, 16#09#),
      835 => to_slv(opcode_type, 16#05#),
      836 => to_slv(opcode_type, 16#0E#),
      837 => to_slv(opcode_type, 16#08#),
      838 => to_slv(opcode_type, 16#10#),
      839 => to_slv(opcode_type, 16#0A#),
      840 => to_slv(opcode_type, 16#09#),
      841 => to_slv(opcode_type, 16#08#),
      842 => to_slv(opcode_type, 16#09#),
      843 => to_slv(opcode_type, 16#0B#),
      844 => to_slv(opcode_type, 16#0F#),
      845 => to_slv(opcode_type, 16#06#),
      846 => to_slv(opcode_type, 16#8C#),
      847 => to_slv(opcode_type, 16#11#),
      848 => to_slv(opcode_type, 16#07#),
      849 => to_slv(opcode_type, 16#09#),
      850 => to_slv(opcode_type, 16#11#),
      851 => to_slv(opcode_type, 16#10#),
      852 => to_slv(opcode_type, 16#08#),
      853 => to_slv(opcode_type, 16#0B#),
      854 => to_slv(opcode_type, 16#0C#),
      855 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#08#),
      865 => to_slv(opcode_type, 16#07#),
      866 => to_slv(opcode_type, 16#01#),
      867 => to_slv(opcode_type, 16#08#),
      868 => to_slv(opcode_type, 16#0D#),
      869 => to_slv(opcode_type, 16#0D#),
      870 => to_slv(opcode_type, 16#09#),
      871 => to_slv(opcode_type, 16#03#),
      872 => to_slv(opcode_type, 16#0C#),
      873 => to_slv(opcode_type, 16#03#),
      874 => to_slv(opcode_type, 16#0A#),
      875 => to_slv(opcode_type, 16#07#),
      876 => to_slv(opcode_type, 16#06#),
      877 => to_slv(opcode_type, 16#03#),
      878 => to_slv(opcode_type, 16#0E#),
      879 => to_slv(opcode_type, 16#01#),
      880 => to_slv(opcode_type, 16#0B#),
      881 => to_slv(opcode_type, 16#06#),
      882 => to_slv(opcode_type, 16#07#),
      883 => to_slv(opcode_type, 16#0B#),
      884 => to_slv(opcode_type, 16#0A#),
      885 => to_slv(opcode_type, 16#03#),
      886 => to_slv(opcode_type, 16#10#),
      887 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#07#),
      898 => to_slv(opcode_type, 16#02#),
      899 => to_slv(opcode_type, 16#07#),
      900 => to_slv(opcode_type, 16#0C#),
      901 => to_slv(opcode_type, 16#0F#),
      902 => to_slv(opcode_type, 16#07#),
      903 => to_slv(opcode_type, 16#07#),
      904 => to_slv(opcode_type, 16#0C#),
      905 => to_slv(opcode_type, 16#0D#),
      906 => to_slv(opcode_type, 16#05#),
      907 => to_slv(opcode_type, 16#0E#),
      908 => to_slv(opcode_type, 16#09#),
      909 => to_slv(opcode_type, 16#01#),
      910 => to_slv(opcode_type, 16#04#),
      911 => to_slv(opcode_type, 16#0E#),
      912 => to_slv(opcode_type, 16#06#),
      913 => to_slv(opcode_type, 16#08#),
      914 => to_slv(opcode_type, 16#0A#),
      915 => to_slv(opcode_type, 16#0D#),
      916 => to_slv(opcode_type, 16#07#),
      917 => to_slv(opcode_type, 16#0C#),
      918 => to_slv(opcode_type, 16#0E#),
      919 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#08#),
      929 => to_slv(opcode_type, 16#02#),
      930 => to_slv(opcode_type, 16#09#),
      931 => to_slv(opcode_type, 16#02#),
      932 => to_slv(opcode_type, 16#0A#),
      933 => to_slv(opcode_type, 16#06#),
      934 => to_slv(opcode_type, 16#0D#),
      935 => to_slv(opcode_type, 16#0E#),
      936 => to_slv(opcode_type, 16#09#),
      937 => to_slv(opcode_type, 16#09#),
      938 => to_slv(opcode_type, 16#07#),
      939 => to_slv(opcode_type, 16#11#),
      940 => to_slv(opcode_type, 16#0F#),
      941 => to_slv(opcode_type, 16#07#),
      942 => to_slv(opcode_type, 16#10#),
      943 => to_slv(opcode_type, 16#0E#),
      944 => to_slv(opcode_type, 16#07#),
      945 => to_slv(opcode_type, 16#09#),
      946 => to_slv(opcode_type, 16#10#),
      947 => to_slv(opcode_type, 16#0B#),
      948 => to_slv(opcode_type, 16#06#),
      949 => to_slv(opcode_type, 16#0C#),
      950 => to_slv(opcode_type, 16#10#),
      951 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#02#),
      962 => to_slv(opcode_type, 16#08#),
      963 => to_slv(opcode_type, 16#02#),
      964 => to_slv(opcode_type, 16#0E#),
      965 => to_slv(opcode_type, 16#08#),
      966 => to_slv(opcode_type, 16#B7#),
      967 => to_slv(opcode_type, 16#11#),
      968 => to_slv(opcode_type, 16#07#),
      969 => to_slv(opcode_type, 16#08#),
      970 => to_slv(opcode_type, 16#09#),
      971 => to_slv(opcode_type, 16#0B#),
      972 => to_slv(opcode_type, 16#0F#),
      973 => to_slv(opcode_type, 16#07#),
      974 => to_slv(opcode_type, 16#0C#),
      975 => to_slv(opcode_type, 16#0D#),
      976 => to_slv(opcode_type, 16#06#),
      977 => to_slv(opcode_type, 16#07#),
      978 => to_slv(opcode_type, 16#0C#),
      979 => to_slv(opcode_type, 16#0A#),
      980 => to_slv(opcode_type, 16#06#),
      981 => to_slv(opcode_type, 16#10#),
      982 => to_slv(opcode_type, 16#0D#),
      983 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#07#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#04#),
      995 => to_slv(opcode_type, 16#05#),
      996 => to_slv(opcode_type, 16#11#),
      997 => to_slv(opcode_type, 16#09#),
      998 => to_slv(opcode_type, 16#06#),
      999 => to_slv(opcode_type, 16#0E#),
      1000 => to_slv(opcode_type, 16#11#),
      1001 => to_slv(opcode_type, 16#04#),
      1002 => to_slv(opcode_type, 16#0F#),
      1003 => to_slv(opcode_type, 16#06#),
      1004 => to_slv(opcode_type, 16#08#),
      1005 => to_slv(opcode_type, 16#09#),
      1006 => to_slv(opcode_type, 16#0C#),
      1007 => to_slv(opcode_type, 16#5D#),
      1008 => to_slv(opcode_type, 16#06#),
      1009 => to_slv(opcode_type, 16#0E#),
      1010 => to_slv(opcode_type, 16#39#),
      1011 => to_slv(opcode_type, 16#01#),
      1012 => to_slv(opcode_type, 16#06#),
      1013 => to_slv(opcode_type, 16#0C#),
      1014 => to_slv(opcode_type, 16#0F#),
      1015 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#06#),
      1025 => to_slv(opcode_type, 16#09#),
      1026 => to_slv(opcode_type, 16#02#),
      1027 => to_slv(opcode_type, 16#04#),
      1028 => to_slv(opcode_type, 16#0D#),
      1029 => to_slv(opcode_type, 16#04#),
      1030 => to_slv(opcode_type, 16#07#),
      1031 => to_slv(opcode_type, 16#0E#),
      1032 => to_slv(opcode_type, 16#0D#),
      1033 => to_slv(opcode_type, 16#06#),
      1034 => to_slv(opcode_type, 16#07#),
      1035 => to_slv(opcode_type, 16#08#),
      1036 => to_slv(opcode_type, 16#0B#),
      1037 => to_slv(opcode_type, 16#0B#),
      1038 => to_slv(opcode_type, 16#09#),
      1039 => to_slv(opcode_type, 16#0C#),
      1040 => to_slv(opcode_type, 16#0C#),
      1041 => to_slv(opcode_type, 16#08#),
      1042 => to_slv(opcode_type, 16#09#),
      1043 => to_slv(opcode_type, 16#0D#),
      1044 => to_slv(opcode_type, 16#0E#),
      1045 => to_slv(opcode_type, 16#03#),
      1046 => to_slv(opcode_type, 16#0D#),
      1047 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#06#),
      1057 => to_slv(opcode_type, 16#03#),
      1058 => to_slv(opcode_type, 16#06#),
      1059 => to_slv(opcode_type, 16#09#),
      1060 => to_slv(opcode_type, 16#0B#),
      1061 => to_slv(opcode_type, 16#0D#),
      1062 => to_slv(opcode_type, 16#08#),
      1063 => to_slv(opcode_type, 16#11#),
      1064 => to_slv(opcode_type, 16#10#),
      1065 => to_slv(opcode_type, 16#09#),
      1066 => to_slv(opcode_type, 16#08#),
      1067 => to_slv(opcode_type, 16#02#),
      1068 => to_slv(opcode_type, 16#90#),
      1069 => to_slv(opcode_type, 16#07#),
      1070 => to_slv(opcode_type, 16#0A#),
      1071 => to_slv(opcode_type, 16#0F#),
      1072 => to_slv(opcode_type, 16#06#),
      1073 => to_slv(opcode_type, 16#08#),
      1074 => to_slv(opcode_type, 16#10#),
      1075 => to_slv(opcode_type, 16#11#),
      1076 => to_slv(opcode_type, 16#06#),
      1077 => to_slv(opcode_type, 16#0A#),
      1078 => to_slv(opcode_type, 16#0C#),
      1079 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#07#),
      1089 => to_slv(opcode_type, 16#02#),
      1090 => to_slv(opcode_type, 16#09#),
      1091 => to_slv(opcode_type, 16#08#),
      1092 => to_slv(opcode_type, 16#11#),
      1093 => to_slv(opcode_type, 16#0E#),
      1094 => to_slv(opcode_type, 16#02#),
      1095 => to_slv(opcode_type, 16#10#),
      1096 => to_slv(opcode_type, 16#07#),
      1097 => to_slv(opcode_type, 16#07#),
      1098 => to_slv(opcode_type, 16#07#),
      1099 => to_slv(opcode_type, 16#0E#),
      1100 => to_slv(opcode_type, 16#0A#),
      1101 => to_slv(opcode_type, 16#08#),
      1102 => to_slv(opcode_type, 16#E3#),
      1103 => to_slv(opcode_type, 16#11#),
      1104 => to_slv(opcode_type, 16#08#),
      1105 => to_slv(opcode_type, 16#06#),
      1106 => to_slv(opcode_type, 16#0E#),
      1107 => to_slv(opcode_type, 16#10#),
      1108 => to_slv(opcode_type, 16#06#),
      1109 => to_slv(opcode_type, 16#11#),
      1110 => to_slv(opcode_type, 16#A2#),
      1111 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#09#),
      1121 => to_slv(opcode_type, 16#07#),
      1122 => to_slv(opcode_type, 16#03#),
      1123 => to_slv(opcode_type, 16#09#),
      1124 => to_slv(opcode_type, 16#0D#),
      1125 => to_slv(opcode_type, 16#0F#),
      1126 => to_slv(opcode_type, 16#02#),
      1127 => to_slv(opcode_type, 16#03#),
      1128 => to_slv(opcode_type, 16#0C#),
      1129 => to_slv(opcode_type, 16#06#),
      1130 => to_slv(opcode_type, 16#07#),
      1131 => to_slv(opcode_type, 16#04#),
      1132 => to_slv(opcode_type, 16#B7#),
      1133 => to_slv(opcode_type, 16#07#),
      1134 => to_slv(opcode_type, 16#0F#),
      1135 => to_slv(opcode_type, 16#0B#),
      1136 => to_slv(opcode_type, 16#08#),
      1137 => to_slv(opcode_type, 16#08#),
      1138 => to_slv(opcode_type, 16#12#),
      1139 => to_slv(opcode_type, 16#11#),
      1140 => to_slv(opcode_type, 16#07#),
      1141 => to_slv(opcode_type, 16#0E#),
      1142 => to_slv(opcode_type, 16#0D#),
      1143 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#09#),
      1153 => to_slv(opcode_type, 16#05#),
      1154 => to_slv(opcode_type, 16#07#),
      1155 => to_slv(opcode_type, 16#01#),
      1156 => to_slv(opcode_type, 16#10#),
      1157 => to_slv(opcode_type, 16#06#),
      1158 => to_slv(opcode_type, 16#40#),
      1159 => to_slv(opcode_type, 16#0F#),
      1160 => to_slv(opcode_type, 16#06#),
      1161 => to_slv(opcode_type, 16#07#),
      1162 => to_slv(opcode_type, 16#07#),
      1163 => to_slv(opcode_type, 16#0C#),
      1164 => to_slv(opcode_type, 16#B0#),
      1165 => to_slv(opcode_type, 16#06#),
      1166 => to_slv(opcode_type, 16#0C#),
      1167 => to_slv(opcode_type, 16#F5#),
      1168 => to_slv(opcode_type, 16#07#),
      1169 => to_slv(opcode_type, 16#06#),
      1170 => to_slv(opcode_type, 16#10#),
      1171 => to_slv(opcode_type, 16#0F#),
      1172 => to_slv(opcode_type, 16#06#),
      1173 => to_slv(opcode_type, 16#11#),
      1174 => to_slv(opcode_type, 16#0D#),
      1175 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#06#),
      1185 => to_slv(opcode_type, 16#07#),
      1186 => to_slv(opcode_type, 16#09#),
      1187 => to_slv(opcode_type, 16#06#),
      1188 => to_slv(opcode_type, 16#0E#),
      1189 => to_slv(opcode_type, 16#10#),
      1190 => to_slv(opcode_type, 16#02#),
      1191 => to_slv(opcode_type, 16#0D#),
      1192 => to_slv(opcode_type, 16#07#),
      1193 => to_slv(opcode_type, 16#03#),
      1194 => to_slv(opcode_type, 16#10#),
      1195 => to_slv(opcode_type, 16#05#),
      1196 => to_slv(opcode_type, 16#0D#),
      1197 => to_slv(opcode_type, 16#06#),
      1198 => to_slv(opcode_type, 16#04#),
      1199 => to_slv(opcode_type, 16#08#),
      1200 => to_slv(opcode_type, 16#0E#),
      1201 => to_slv(opcode_type, 16#0E#),
      1202 => to_slv(opcode_type, 16#08#),
      1203 => to_slv(opcode_type, 16#07#),
      1204 => to_slv(opcode_type, 16#0E#),
      1205 => to_slv(opcode_type, 16#0B#),
      1206 => to_slv(opcode_type, 16#11#),
      1207 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#09#),
      1217 => to_slv(opcode_type, 16#07#),
      1218 => to_slv(opcode_type, 16#04#),
      1219 => to_slv(opcode_type, 16#06#),
      1220 => to_slv(opcode_type, 16#0F#),
      1221 => to_slv(opcode_type, 16#10#),
      1222 => to_slv(opcode_type, 16#05#),
      1223 => to_slv(opcode_type, 16#03#),
      1224 => to_slv(opcode_type, 16#11#),
      1225 => to_slv(opcode_type, 16#06#),
      1226 => to_slv(opcode_type, 16#09#),
      1227 => to_slv(opcode_type, 16#06#),
      1228 => to_slv(opcode_type, 16#0C#),
      1229 => to_slv(opcode_type, 16#11#),
      1230 => to_slv(opcode_type, 16#01#),
      1231 => to_slv(opcode_type, 16#11#),
      1232 => to_slv(opcode_type, 16#06#),
      1233 => to_slv(opcode_type, 16#08#),
      1234 => to_slv(opcode_type, 16#0C#),
      1235 => to_slv(opcode_type, 16#0C#),
      1236 => to_slv(opcode_type, 16#08#),
      1237 => to_slv(opcode_type, 16#73#),
      1238 => to_slv(opcode_type, 16#0F#),
      1239 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#09#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#07#),
      1251 => to_slv(opcode_type, 16#05#),
      1252 => to_slv(opcode_type, 16#0F#),
      1253 => to_slv(opcode_type, 16#03#),
      1254 => to_slv(opcode_type, 16#10#),
      1255 => to_slv(opcode_type, 16#07#),
      1256 => to_slv(opcode_type, 16#05#),
      1257 => to_slv(opcode_type, 16#10#),
      1258 => to_slv(opcode_type, 16#09#),
      1259 => to_slv(opcode_type, 16#0B#),
      1260 => to_slv(opcode_type, 16#0B#),
      1261 => to_slv(opcode_type, 16#09#),
      1262 => to_slv(opcode_type, 16#07#),
      1263 => to_slv(opcode_type, 16#09#),
      1264 => to_slv(opcode_type, 16#0D#),
      1265 => to_slv(opcode_type, 16#0B#),
      1266 => to_slv(opcode_type, 16#01#),
      1267 => to_slv(opcode_type, 16#0A#),
      1268 => to_slv(opcode_type, 16#08#),
      1269 => to_slv(opcode_type, 16#0C#),
      1270 => to_slv(opcode_type, 16#7E#),
      1271 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#08#),
      1281 => to_slv(opcode_type, 16#05#),
      1282 => to_slv(opcode_type, 16#09#),
      1283 => to_slv(opcode_type, 16#03#),
      1284 => to_slv(opcode_type, 16#0B#),
      1285 => to_slv(opcode_type, 16#06#),
      1286 => to_slv(opcode_type, 16#0B#),
      1287 => to_slv(opcode_type, 16#0F#),
      1288 => to_slv(opcode_type, 16#06#),
      1289 => to_slv(opcode_type, 16#08#),
      1290 => to_slv(opcode_type, 16#06#),
      1291 => to_slv(opcode_type, 16#0E#),
      1292 => to_slv(opcode_type, 16#0C#),
      1293 => to_slv(opcode_type, 16#09#),
      1294 => to_slv(opcode_type, 16#0F#),
      1295 => to_slv(opcode_type, 16#0E#),
      1296 => to_slv(opcode_type, 16#09#),
      1297 => to_slv(opcode_type, 16#09#),
      1298 => to_slv(opcode_type, 16#0A#),
      1299 => to_slv(opcode_type, 16#0E#),
      1300 => to_slv(opcode_type, 16#08#),
      1301 => to_slv(opcode_type, 16#0D#),
      1302 => to_slv(opcode_type, 16#55#),
      1303 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#06#),
      1313 => to_slv(opcode_type, 16#02#),
      1314 => to_slv(opcode_type, 16#09#),
      1315 => to_slv(opcode_type, 16#09#),
      1316 => to_slv(opcode_type, 16#0E#),
      1317 => to_slv(opcode_type, 16#0B#),
      1318 => to_slv(opcode_type, 16#05#),
      1319 => to_slv(opcode_type, 16#0F#),
      1320 => to_slv(opcode_type, 16#09#),
      1321 => to_slv(opcode_type, 16#08#),
      1322 => to_slv(opcode_type, 16#09#),
      1323 => to_slv(opcode_type, 16#0E#),
      1324 => to_slv(opcode_type, 16#C4#),
      1325 => to_slv(opcode_type, 16#07#),
      1326 => to_slv(opcode_type, 16#37#),
      1327 => to_slv(opcode_type, 16#11#),
      1328 => to_slv(opcode_type, 16#07#),
      1329 => to_slv(opcode_type, 16#09#),
      1330 => to_slv(opcode_type, 16#0A#),
      1331 => to_slv(opcode_type, 16#11#),
      1332 => to_slv(opcode_type, 16#08#),
      1333 => to_slv(opcode_type, 16#0C#),
      1334 => to_slv(opcode_type, 16#0D#),
      1335 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#09#),
      1345 => to_slv(opcode_type, 16#07#),
      1346 => to_slv(opcode_type, 16#09#),
      1347 => to_slv(opcode_type, 16#03#),
      1348 => to_slv(opcode_type, 16#0E#),
      1349 => to_slv(opcode_type, 16#09#),
      1350 => to_slv(opcode_type, 16#10#),
      1351 => to_slv(opcode_type, 16#0D#),
      1352 => to_slv(opcode_type, 16#02#),
      1353 => to_slv(opcode_type, 16#09#),
      1354 => to_slv(opcode_type, 16#0C#),
      1355 => to_slv(opcode_type, 16#11#),
      1356 => to_slv(opcode_type, 16#07#),
      1357 => to_slv(opcode_type, 16#07#),
      1358 => to_slv(opcode_type, 16#09#),
      1359 => to_slv(opcode_type, 16#0E#),
      1360 => to_slv(opcode_type, 16#11#),
      1361 => to_slv(opcode_type, 16#06#),
      1362 => to_slv(opcode_type, 16#0C#),
      1363 => to_slv(opcode_type, 16#11#),
      1364 => to_slv(opcode_type, 16#08#),
      1365 => to_slv(opcode_type, 16#0C#),
      1366 => to_slv(opcode_type, 16#0F#),
      1367 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#07#),
      1377 => to_slv(opcode_type, 16#06#),
      1378 => to_slv(opcode_type, 16#01#),
      1379 => to_slv(opcode_type, 16#08#),
      1380 => to_slv(opcode_type, 16#0A#),
      1381 => to_slv(opcode_type, 16#0C#),
      1382 => to_slv(opcode_type, 16#06#),
      1383 => to_slv(opcode_type, 16#09#),
      1384 => to_slv(opcode_type, 16#0E#),
      1385 => to_slv(opcode_type, 16#0A#),
      1386 => to_slv(opcode_type, 16#05#),
      1387 => to_slv(opcode_type, 16#0D#),
      1388 => to_slv(opcode_type, 16#08#),
      1389 => to_slv(opcode_type, 16#05#),
      1390 => to_slv(opcode_type, 16#03#),
      1391 => to_slv(opcode_type, 16#0A#),
      1392 => to_slv(opcode_type, 16#06#),
      1393 => to_slv(opcode_type, 16#06#),
      1394 => to_slv(opcode_type, 16#0C#),
      1395 => to_slv(opcode_type, 16#0A#),
      1396 => to_slv(opcode_type, 16#06#),
      1397 => to_slv(opcode_type, 16#A7#),
      1398 => to_slv(opcode_type, 16#11#),
      1399 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#08#),
      1410 => to_slv(opcode_type, 16#05#),
      1411 => to_slv(opcode_type, 16#06#),
      1412 => to_slv(opcode_type, 16#0E#),
      1413 => to_slv(opcode_type, 16#0D#),
      1414 => to_slv(opcode_type, 16#09#),
      1415 => to_slv(opcode_type, 16#03#),
      1416 => to_slv(opcode_type, 16#0A#),
      1417 => to_slv(opcode_type, 16#04#),
      1418 => to_slv(opcode_type, 16#F5#),
      1419 => to_slv(opcode_type, 16#09#),
      1420 => to_slv(opcode_type, 16#01#),
      1421 => to_slv(opcode_type, 16#09#),
      1422 => to_slv(opcode_type, 16#10#),
      1423 => to_slv(opcode_type, 16#0A#),
      1424 => to_slv(opcode_type, 16#07#),
      1425 => to_slv(opcode_type, 16#06#),
      1426 => to_slv(opcode_type, 16#0C#),
      1427 => to_slv(opcode_type, 16#0F#),
      1428 => to_slv(opcode_type, 16#08#),
      1429 => to_slv(opcode_type, 16#0C#),
      1430 => to_slv(opcode_type, 16#0F#),
      1431 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#09#),
      1441 => to_slv(opcode_type, 16#02#),
      1442 => to_slv(opcode_type, 16#06#),
      1443 => to_slv(opcode_type, 16#04#),
      1444 => to_slv(opcode_type, 16#E7#),
      1445 => to_slv(opcode_type, 16#08#),
      1446 => to_slv(opcode_type, 16#0F#),
      1447 => to_slv(opcode_type, 16#11#),
      1448 => to_slv(opcode_type, 16#07#),
      1449 => to_slv(opcode_type, 16#09#),
      1450 => to_slv(opcode_type, 16#08#),
      1451 => to_slv(opcode_type, 16#0A#),
      1452 => to_slv(opcode_type, 16#0A#),
      1453 => to_slv(opcode_type, 16#07#),
      1454 => to_slv(opcode_type, 16#0E#),
      1455 => to_slv(opcode_type, 16#0D#),
      1456 => to_slv(opcode_type, 16#06#),
      1457 => to_slv(opcode_type, 16#06#),
      1458 => to_slv(opcode_type, 16#0B#),
      1459 => to_slv(opcode_type, 16#0F#),
      1460 => to_slv(opcode_type, 16#08#),
      1461 => to_slv(opcode_type, 16#0E#),
      1462 => to_slv(opcode_type, 16#11#),
      1463 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#08#),
      1473 => to_slv(opcode_type, 16#02#),
      1474 => to_slv(opcode_type, 16#07#),
      1475 => to_slv(opcode_type, 16#04#),
      1476 => to_slv(opcode_type, 16#0A#),
      1477 => to_slv(opcode_type, 16#06#),
      1478 => to_slv(opcode_type, 16#11#),
      1479 => to_slv(opcode_type, 16#22#),
      1480 => to_slv(opcode_type, 16#08#),
      1481 => to_slv(opcode_type, 16#07#),
      1482 => to_slv(opcode_type, 16#09#),
      1483 => to_slv(opcode_type, 16#0F#),
      1484 => to_slv(opcode_type, 16#0E#),
      1485 => to_slv(opcode_type, 16#07#),
      1486 => to_slv(opcode_type, 16#0B#),
      1487 => to_slv(opcode_type, 16#0C#),
      1488 => to_slv(opcode_type, 16#08#),
      1489 => to_slv(opcode_type, 16#07#),
      1490 => to_slv(opcode_type, 16#8C#),
      1491 => to_slv(opcode_type, 16#0B#),
      1492 => to_slv(opcode_type, 16#09#),
      1493 => to_slv(opcode_type, 16#0F#),
      1494 => to_slv(opcode_type, 16#0A#),
      1495 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#07#),
      1505 => to_slv(opcode_type, 16#06#),
      1506 => to_slv(opcode_type, 16#05#),
      1507 => to_slv(opcode_type, 16#05#),
      1508 => to_slv(opcode_type, 16#0B#),
      1509 => to_slv(opcode_type, 16#07#),
      1510 => to_slv(opcode_type, 16#05#),
      1511 => to_slv(opcode_type, 16#0B#),
      1512 => to_slv(opcode_type, 16#04#),
      1513 => to_slv(opcode_type, 16#0F#),
      1514 => to_slv(opcode_type, 16#08#),
      1515 => to_slv(opcode_type, 16#09#),
      1516 => to_slv(opcode_type, 16#04#),
      1517 => to_slv(opcode_type, 16#11#),
      1518 => to_slv(opcode_type, 16#06#),
      1519 => to_slv(opcode_type, 16#58#),
      1520 => to_slv(opcode_type, 16#0C#),
      1521 => to_slv(opcode_type, 16#07#),
      1522 => to_slv(opcode_type, 16#02#),
      1523 => to_slv(opcode_type, 16#0C#),
      1524 => to_slv(opcode_type, 16#07#),
      1525 => to_slv(opcode_type, 16#11#),
      1526 => to_slv(opcode_type, 16#0F#),
      1527 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#08#),
      1537 => to_slv(opcode_type, 16#01#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#03#),
      1540 => to_slv(opcode_type, 16#0E#),
      1541 => to_slv(opcode_type, 16#08#),
      1542 => to_slv(opcode_type, 16#0C#),
      1543 => to_slv(opcode_type, 16#11#),
      1544 => to_slv(opcode_type, 16#06#),
      1545 => to_slv(opcode_type, 16#06#),
      1546 => to_slv(opcode_type, 16#07#),
      1547 => to_slv(opcode_type, 16#10#),
      1548 => to_slv(opcode_type, 16#0A#),
      1549 => to_slv(opcode_type, 16#09#),
      1550 => to_slv(opcode_type, 16#0C#),
      1551 => to_slv(opcode_type, 16#10#),
      1552 => to_slv(opcode_type, 16#06#),
      1553 => to_slv(opcode_type, 16#07#),
      1554 => to_slv(opcode_type, 16#5A#),
      1555 => to_slv(opcode_type, 16#0C#),
      1556 => to_slv(opcode_type, 16#09#),
      1557 => to_slv(opcode_type, 16#0E#),
      1558 => to_slv(opcode_type, 16#0B#),
      1559 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#06#),
      1569 => to_slv(opcode_type, 16#09#),
      1570 => to_slv(opcode_type, 16#08#),
      1571 => to_slv(opcode_type, 16#05#),
      1572 => to_slv(opcode_type, 16#0F#),
      1573 => to_slv(opcode_type, 16#08#),
      1574 => to_slv(opcode_type, 16#0B#),
      1575 => to_slv(opcode_type, 16#0E#),
      1576 => to_slv(opcode_type, 16#02#),
      1577 => to_slv(opcode_type, 16#07#),
      1578 => to_slv(opcode_type, 16#10#),
      1579 => to_slv(opcode_type, 16#10#),
      1580 => to_slv(opcode_type, 16#09#),
      1581 => to_slv(opcode_type, 16#03#),
      1582 => to_slv(opcode_type, 16#05#),
      1583 => to_slv(opcode_type, 16#F9#),
      1584 => to_slv(opcode_type, 16#08#),
      1585 => to_slv(opcode_type, 16#07#),
      1586 => to_slv(opcode_type, 16#0F#),
      1587 => to_slv(opcode_type, 16#0E#),
      1588 => to_slv(opcode_type, 16#06#),
      1589 => to_slv(opcode_type, 16#4F#),
      1590 => to_slv(opcode_type, 16#10#),
      1591 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#08#),
      1601 => to_slv(opcode_type, 16#07#),
      1602 => to_slv(opcode_type, 16#04#),
      1603 => to_slv(opcode_type, 16#02#),
      1604 => to_slv(opcode_type, 16#11#),
      1605 => to_slv(opcode_type, 16#03#),
      1606 => to_slv(opcode_type, 16#08#),
      1607 => to_slv(opcode_type, 16#10#),
      1608 => to_slv(opcode_type, 16#0B#),
      1609 => to_slv(opcode_type, 16#07#),
      1610 => to_slv(opcode_type, 16#06#),
      1611 => to_slv(opcode_type, 16#04#),
      1612 => to_slv(opcode_type, 16#0B#),
      1613 => to_slv(opcode_type, 16#07#),
      1614 => to_slv(opcode_type, 16#0B#),
      1615 => to_slv(opcode_type, 16#0D#),
      1616 => to_slv(opcode_type, 16#07#),
      1617 => to_slv(opcode_type, 16#06#),
      1618 => to_slv(opcode_type, 16#0C#),
      1619 => to_slv(opcode_type, 16#0E#),
      1620 => to_slv(opcode_type, 16#06#),
      1621 => to_slv(opcode_type, 16#0F#),
      1622 => to_slv(opcode_type, 16#0F#),
      1623 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#07#),
      1633 => to_slv(opcode_type, 16#09#),
      1634 => to_slv(opcode_type, 16#06#),
      1635 => to_slv(opcode_type, 16#04#),
      1636 => to_slv(opcode_type, 16#0F#),
      1637 => to_slv(opcode_type, 16#01#),
      1638 => to_slv(opcode_type, 16#0E#),
      1639 => to_slv(opcode_type, 16#07#),
      1640 => to_slv(opcode_type, 16#01#),
      1641 => to_slv(opcode_type, 16#0C#),
      1642 => to_slv(opcode_type, 16#08#),
      1643 => to_slv(opcode_type, 16#0B#),
      1644 => to_slv(opcode_type, 16#0E#),
      1645 => to_slv(opcode_type, 16#06#),
      1646 => to_slv(opcode_type, 16#04#),
      1647 => to_slv(opcode_type, 16#06#),
      1648 => to_slv(opcode_type, 16#0D#),
      1649 => to_slv(opcode_type, 16#0B#),
      1650 => to_slv(opcode_type, 16#06#),
      1651 => to_slv(opcode_type, 16#09#),
      1652 => to_slv(opcode_type, 16#11#),
      1653 => to_slv(opcode_type, 16#10#),
      1654 => to_slv(opcode_type, 16#11#),
      1655 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#05#),
      1666 => to_slv(opcode_type, 16#06#),
      1667 => to_slv(opcode_type, 16#09#),
      1668 => to_slv(opcode_type, 16#0D#),
      1669 => to_slv(opcode_type, 16#0D#),
      1670 => to_slv(opcode_type, 16#03#),
      1671 => to_slv(opcode_type, 16#0E#),
      1672 => to_slv(opcode_type, 16#06#),
      1673 => to_slv(opcode_type, 16#08#),
      1674 => to_slv(opcode_type, 16#06#),
      1675 => to_slv(opcode_type, 16#85#),
      1676 => to_slv(opcode_type, 16#0C#),
      1677 => to_slv(opcode_type, 16#06#),
      1678 => to_slv(opcode_type, 16#0D#),
      1679 => to_slv(opcode_type, 16#10#),
      1680 => to_slv(opcode_type, 16#06#),
      1681 => to_slv(opcode_type, 16#07#),
      1682 => to_slv(opcode_type, 16#0D#),
      1683 => to_slv(opcode_type, 16#0D#),
      1684 => to_slv(opcode_type, 16#06#),
      1685 => to_slv(opcode_type, 16#11#),
      1686 => to_slv(opcode_type, 16#0D#),
      1687 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#09#),
      1697 => to_slv(opcode_type, 16#02#),
      1698 => to_slv(opcode_type, 16#06#),
      1699 => to_slv(opcode_type, 16#04#),
      1700 => to_slv(opcode_type, 16#0D#),
      1701 => to_slv(opcode_type, 16#09#),
      1702 => to_slv(opcode_type, 16#0F#),
      1703 => to_slv(opcode_type, 16#0F#),
      1704 => to_slv(opcode_type, 16#09#),
      1705 => to_slv(opcode_type, 16#06#),
      1706 => to_slv(opcode_type, 16#08#),
      1707 => to_slv(opcode_type, 16#0A#),
      1708 => to_slv(opcode_type, 16#11#),
      1709 => to_slv(opcode_type, 16#07#),
      1710 => to_slv(opcode_type, 16#10#),
      1711 => to_slv(opcode_type, 16#10#),
      1712 => to_slv(opcode_type, 16#07#),
      1713 => to_slv(opcode_type, 16#06#),
      1714 => to_slv(opcode_type, 16#0D#),
      1715 => to_slv(opcode_type, 16#0E#),
      1716 => to_slv(opcode_type, 16#09#),
      1717 => to_slv(opcode_type, 16#0E#),
      1718 => to_slv(opcode_type, 16#0F#),
      1719 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#06#),
      1729 => to_slv(opcode_type, 16#02#),
      1730 => to_slv(opcode_type, 16#09#),
      1731 => to_slv(opcode_type, 16#04#),
      1732 => to_slv(opcode_type, 16#0C#),
      1733 => to_slv(opcode_type, 16#09#),
      1734 => to_slv(opcode_type, 16#0D#),
      1735 => to_slv(opcode_type, 16#0C#),
      1736 => to_slv(opcode_type, 16#07#),
      1737 => to_slv(opcode_type, 16#09#),
      1738 => to_slv(opcode_type, 16#07#),
      1739 => to_slv(opcode_type, 16#0C#),
      1740 => to_slv(opcode_type, 16#0F#),
      1741 => to_slv(opcode_type, 16#07#),
      1742 => to_slv(opcode_type, 16#0A#),
      1743 => to_slv(opcode_type, 16#0A#),
      1744 => to_slv(opcode_type, 16#06#),
      1745 => to_slv(opcode_type, 16#07#),
      1746 => to_slv(opcode_type, 16#0D#),
      1747 => to_slv(opcode_type, 16#DB#),
      1748 => to_slv(opcode_type, 16#08#),
      1749 => to_slv(opcode_type, 16#0A#),
      1750 => to_slv(opcode_type, 16#0D#),
      1751 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#07#),
      1761 => to_slv(opcode_type, 16#02#),
      1762 => to_slv(opcode_type, 16#07#),
      1763 => to_slv(opcode_type, 16#09#),
      1764 => to_slv(opcode_type, 16#0C#),
      1765 => to_slv(opcode_type, 16#0B#),
      1766 => to_slv(opcode_type, 16#06#),
      1767 => to_slv(opcode_type, 16#0D#),
      1768 => to_slv(opcode_type, 16#EB#),
      1769 => to_slv(opcode_type, 16#08#),
      1770 => to_slv(opcode_type, 16#09#),
      1771 => to_slv(opcode_type, 16#01#),
      1772 => to_slv(opcode_type, 16#0D#),
      1773 => to_slv(opcode_type, 16#09#),
      1774 => to_slv(opcode_type, 16#10#),
      1775 => to_slv(opcode_type, 16#0D#),
      1776 => to_slv(opcode_type, 16#07#),
      1777 => to_slv(opcode_type, 16#07#),
      1778 => to_slv(opcode_type, 16#0C#),
      1779 => to_slv(opcode_type, 16#0B#),
      1780 => to_slv(opcode_type, 16#07#),
      1781 => to_slv(opcode_type, 16#0B#),
      1782 => to_slv(opcode_type, 16#0C#),
      1783 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#09#),
      1793 => to_slv(opcode_type, 16#04#),
      1794 => to_slv(opcode_type, 16#06#),
      1795 => to_slv(opcode_type, 16#07#),
      1796 => to_slv(opcode_type, 16#0B#),
      1797 => to_slv(opcode_type, 16#10#),
      1798 => to_slv(opcode_type, 16#01#),
      1799 => to_slv(opcode_type, 16#0F#),
      1800 => to_slv(opcode_type, 16#09#),
      1801 => to_slv(opcode_type, 16#07#),
      1802 => to_slv(opcode_type, 16#09#),
      1803 => to_slv(opcode_type, 16#10#),
      1804 => to_slv(opcode_type, 16#0B#),
      1805 => to_slv(opcode_type, 16#09#),
      1806 => to_slv(opcode_type, 16#11#),
      1807 => to_slv(opcode_type, 16#0B#),
      1808 => to_slv(opcode_type, 16#09#),
      1809 => to_slv(opcode_type, 16#06#),
      1810 => to_slv(opcode_type, 16#0F#),
      1811 => to_slv(opcode_type, 16#10#),
      1812 => to_slv(opcode_type, 16#07#),
      1813 => to_slv(opcode_type, 16#0D#),
      1814 => to_slv(opcode_type, 16#27#),
      1815 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#09#),
      1825 => to_slv(opcode_type, 16#08#),
      1826 => to_slv(opcode_type, 16#08#),
      1827 => to_slv(opcode_type, 16#05#),
      1828 => to_slv(opcode_type, 16#0E#),
      1829 => to_slv(opcode_type, 16#09#),
      1830 => to_slv(opcode_type, 16#0F#),
      1831 => to_slv(opcode_type, 16#0C#),
      1832 => to_slv(opcode_type, 16#09#),
      1833 => to_slv(opcode_type, 16#04#),
      1834 => to_slv(opcode_type, 16#0E#),
      1835 => to_slv(opcode_type, 16#09#),
      1836 => to_slv(opcode_type, 16#0D#),
      1837 => to_slv(opcode_type, 16#0D#),
      1838 => to_slv(opcode_type, 16#07#),
      1839 => to_slv(opcode_type, 16#02#),
      1840 => to_slv(opcode_type, 16#04#),
      1841 => to_slv(opcode_type, 16#0F#),
      1842 => to_slv(opcode_type, 16#08#),
      1843 => to_slv(opcode_type, 16#06#),
      1844 => to_slv(opcode_type, 16#0C#),
      1845 => to_slv(opcode_type, 16#11#),
      1846 => to_slv(opcode_type, 16#E9#),
      1847 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#06#),
      1857 => to_slv(opcode_type, 16#09#),
      1858 => to_slv(opcode_type, 16#07#),
      1859 => to_slv(opcode_type, 16#09#),
      1860 => to_slv(opcode_type, 16#0F#),
      1861 => to_slv(opcode_type, 16#F5#),
      1862 => to_slv(opcode_type, 16#06#),
      1863 => to_slv(opcode_type, 16#0C#),
      1864 => to_slv(opcode_type, 16#0A#),
      1865 => to_slv(opcode_type, 16#07#),
      1866 => to_slv(opcode_type, 16#02#),
      1867 => to_slv(opcode_type, 16#0E#),
      1868 => to_slv(opcode_type, 16#01#),
      1869 => to_slv(opcode_type, 16#0A#),
      1870 => to_slv(opcode_type, 16#06#),
      1871 => to_slv(opcode_type, 16#02#),
      1872 => to_slv(opcode_type, 16#04#),
      1873 => to_slv(opcode_type, 16#0C#),
      1874 => to_slv(opcode_type, 16#07#),
      1875 => to_slv(opcode_type, 16#06#),
      1876 => to_slv(opcode_type, 16#0C#),
      1877 => to_slv(opcode_type, 16#11#),
      1878 => to_slv(opcode_type, 16#11#),
      1879 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#07#),
      1890 => to_slv(opcode_type, 16#02#),
      1891 => to_slv(opcode_type, 16#03#),
      1892 => to_slv(opcode_type, 16#11#),
      1893 => to_slv(opcode_type, 16#01#),
      1894 => to_slv(opcode_type, 16#03#),
      1895 => to_slv(opcode_type, 16#0A#),
      1896 => to_slv(opcode_type, 16#09#),
      1897 => to_slv(opcode_type, 16#07#),
      1898 => to_slv(opcode_type, 16#09#),
      1899 => to_slv(opcode_type, 16#11#),
      1900 => to_slv(opcode_type, 16#0C#),
      1901 => to_slv(opcode_type, 16#06#),
      1902 => to_slv(opcode_type, 16#0F#),
      1903 => to_slv(opcode_type, 16#0D#),
      1904 => to_slv(opcode_type, 16#07#),
      1905 => to_slv(opcode_type, 16#09#),
      1906 => to_slv(opcode_type, 16#3A#),
      1907 => to_slv(opcode_type, 16#0C#),
      1908 => to_slv(opcode_type, 16#06#),
      1909 => to_slv(opcode_type, 16#FC#),
      1910 => to_slv(opcode_type, 16#0C#),
      1911 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#08#),
      1921 => to_slv(opcode_type, 16#08#),
      1922 => to_slv(opcode_type, 16#02#),
      1923 => to_slv(opcode_type, 16#08#),
      1924 => to_slv(opcode_type, 16#0C#),
      1925 => to_slv(opcode_type, 16#0F#),
      1926 => to_slv(opcode_type, 16#08#),
      1927 => to_slv(opcode_type, 16#01#),
      1928 => to_slv(opcode_type, 16#0F#),
      1929 => to_slv(opcode_type, 16#04#),
      1930 => to_slv(opcode_type, 16#0A#),
      1931 => to_slv(opcode_type, 16#06#),
      1932 => to_slv(opcode_type, 16#05#),
      1933 => to_slv(opcode_type, 16#07#),
      1934 => to_slv(opcode_type, 16#0D#),
      1935 => to_slv(opcode_type, 16#10#),
      1936 => to_slv(opcode_type, 16#06#),
      1937 => to_slv(opcode_type, 16#08#),
      1938 => to_slv(opcode_type, 16#0F#),
      1939 => to_slv(opcode_type, 16#11#),
      1940 => to_slv(opcode_type, 16#09#),
      1941 => to_slv(opcode_type, 16#0C#),
      1942 => to_slv(opcode_type, 16#0A#),
      1943 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#07#),
      1953 => to_slv(opcode_type, 16#06#),
      1954 => to_slv(opcode_type, 16#08#),
      1955 => to_slv(opcode_type, 16#03#),
      1956 => to_slv(opcode_type, 16#0A#),
      1957 => to_slv(opcode_type, 16#04#),
      1958 => to_slv(opcode_type, 16#0C#),
      1959 => to_slv(opcode_type, 16#06#),
      1960 => to_slv(opcode_type, 16#02#),
      1961 => to_slv(opcode_type, 16#11#),
      1962 => to_slv(opcode_type, 16#09#),
      1963 => to_slv(opcode_type, 16#0A#),
      1964 => to_slv(opcode_type, 16#11#),
      1965 => to_slv(opcode_type, 16#06#),
      1966 => to_slv(opcode_type, 16#08#),
      1967 => to_slv(opcode_type, 16#01#),
      1968 => to_slv(opcode_type, 16#0E#),
      1969 => to_slv(opcode_type, 16#09#),
      1970 => to_slv(opcode_type, 16#11#),
      1971 => to_slv(opcode_type, 16#0D#),
      1972 => to_slv(opcode_type, 16#07#),
      1973 => to_slv(opcode_type, 16#0E#),
      1974 => to_slv(opcode_type, 16#0D#),
      1975 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#08#),
      1985 => to_slv(opcode_type, 16#05#),
      1986 => to_slv(opcode_type, 16#07#),
      1987 => to_slv(opcode_type, 16#02#),
      1988 => to_slv(opcode_type, 16#0C#),
      1989 => to_slv(opcode_type, 16#08#),
      1990 => to_slv(opcode_type, 16#0F#),
      1991 => to_slv(opcode_type, 16#38#),
      1992 => to_slv(opcode_type, 16#09#),
      1993 => to_slv(opcode_type, 16#08#),
      1994 => to_slv(opcode_type, 16#06#),
      1995 => to_slv(opcode_type, 16#0B#),
      1996 => to_slv(opcode_type, 16#0C#),
      1997 => to_slv(opcode_type, 16#08#),
      1998 => to_slv(opcode_type, 16#C2#),
      1999 => to_slv(opcode_type, 16#0F#),
      2000 => to_slv(opcode_type, 16#06#),
      2001 => to_slv(opcode_type, 16#09#),
      2002 => to_slv(opcode_type, 16#0F#),
      2003 => to_slv(opcode_type, 16#0B#),
      2004 => to_slv(opcode_type, 16#08#),
      2005 => to_slv(opcode_type, 16#B0#),
      2006 => to_slv(opcode_type, 16#0A#),
      2007 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#08#),
      2017 => to_slv(opcode_type, 16#04#),
      2018 => to_slv(opcode_type, 16#06#),
      2019 => to_slv(opcode_type, 16#05#),
      2020 => to_slv(opcode_type, 16#0F#),
      2021 => to_slv(opcode_type, 16#07#),
      2022 => to_slv(opcode_type, 16#10#),
      2023 => to_slv(opcode_type, 16#11#),
      2024 => to_slv(opcode_type, 16#07#),
      2025 => to_slv(opcode_type, 16#06#),
      2026 => to_slv(opcode_type, 16#09#),
      2027 => to_slv(opcode_type, 16#0C#),
      2028 => to_slv(opcode_type, 16#0F#),
      2029 => to_slv(opcode_type, 16#09#),
      2030 => to_slv(opcode_type, 16#0E#),
      2031 => to_slv(opcode_type, 16#0C#),
      2032 => to_slv(opcode_type, 16#09#),
      2033 => to_slv(opcode_type, 16#06#),
      2034 => to_slv(opcode_type, 16#11#),
      2035 => to_slv(opcode_type, 16#0C#),
      2036 => to_slv(opcode_type, 16#07#),
      2037 => to_slv(opcode_type, 16#0D#),
      2038 => to_slv(opcode_type, 16#11#),
      2039 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#09#),
      2049 => to_slv(opcode_type, 16#07#),
      2050 => to_slv(opcode_type, 16#07#),
      2051 => to_slv(opcode_type, 16#08#),
      2052 => to_slv(opcode_type, 16#0F#),
      2053 => to_slv(opcode_type, 16#0C#),
      2054 => to_slv(opcode_type, 16#01#),
      2055 => to_slv(opcode_type, 16#0C#),
      2056 => to_slv(opcode_type, 16#03#),
      2057 => to_slv(opcode_type, 16#02#),
      2058 => to_slv(opcode_type, 16#0D#),
      2059 => to_slv(opcode_type, 16#09#),
      2060 => to_slv(opcode_type, 16#06#),
      2061 => to_slv(opcode_type, 16#02#),
      2062 => to_slv(opcode_type, 16#0A#),
      2063 => to_slv(opcode_type, 16#08#),
      2064 => to_slv(opcode_type, 16#0B#),
      2065 => to_slv(opcode_type, 16#0B#),
      2066 => to_slv(opcode_type, 16#07#),
      2067 => to_slv(opcode_type, 16#03#),
      2068 => to_slv(opcode_type, 16#0F#),
      2069 => to_slv(opcode_type, 16#05#),
      2070 => to_slv(opcode_type, 16#0C#),
      2071 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#08#),
      2081 => to_slv(opcode_type, 16#04#),
      2082 => to_slv(opcode_type, 16#08#),
      2083 => to_slv(opcode_type, 16#01#),
      2084 => to_slv(opcode_type, 16#0F#),
      2085 => to_slv(opcode_type, 16#07#),
      2086 => to_slv(opcode_type, 16#DB#),
      2087 => to_slv(opcode_type, 16#0C#),
      2088 => to_slv(opcode_type, 16#08#),
      2089 => to_slv(opcode_type, 16#09#),
      2090 => to_slv(opcode_type, 16#08#),
      2091 => to_slv(opcode_type, 16#0B#),
      2092 => to_slv(opcode_type, 16#0E#),
      2093 => to_slv(opcode_type, 16#08#),
      2094 => to_slv(opcode_type, 16#10#),
      2095 => to_slv(opcode_type, 16#0E#),
      2096 => to_slv(opcode_type, 16#09#),
      2097 => to_slv(opcode_type, 16#06#),
      2098 => to_slv(opcode_type, 16#0F#),
      2099 => to_slv(opcode_type, 16#11#),
      2100 => to_slv(opcode_type, 16#09#),
      2101 => to_slv(opcode_type, 16#0B#),
      2102 => to_slv(opcode_type, 16#0E#),
      2103 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#08#),
      2113 => to_slv(opcode_type, 16#02#),
      2114 => to_slv(opcode_type, 16#08#),
      2115 => to_slv(opcode_type, 16#09#),
      2116 => to_slv(opcode_type, 16#0E#),
      2117 => to_slv(opcode_type, 16#D5#),
      2118 => to_slv(opcode_type, 16#08#),
      2119 => to_slv(opcode_type, 16#0A#),
      2120 => to_slv(opcode_type, 16#0A#),
      2121 => to_slv(opcode_type, 16#07#),
      2122 => to_slv(opcode_type, 16#08#),
      2123 => to_slv(opcode_type, 16#03#),
      2124 => to_slv(opcode_type, 16#0C#),
      2125 => to_slv(opcode_type, 16#09#),
      2126 => to_slv(opcode_type, 16#10#),
      2127 => to_slv(opcode_type, 16#0B#),
      2128 => to_slv(opcode_type, 16#09#),
      2129 => to_slv(opcode_type, 16#09#),
      2130 => to_slv(opcode_type, 16#11#),
      2131 => to_slv(opcode_type, 16#0F#),
      2132 => to_slv(opcode_type, 16#09#),
      2133 => to_slv(opcode_type, 16#0E#),
      2134 => to_slv(opcode_type, 16#0A#),
      2135 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#09#),
      2146 => to_slv(opcode_type, 16#09#),
      2147 => to_slv(opcode_type, 16#05#),
      2148 => to_slv(opcode_type, 16#11#),
      2149 => to_slv(opcode_type, 16#08#),
      2150 => to_slv(opcode_type, 16#0D#),
      2151 => to_slv(opcode_type, 16#0D#),
      2152 => to_slv(opcode_type, 16#01#),
      2153 => to_slv(opcode_type, 16#05#),
      2154 => to_slv(opcode_type, 16#0A#),
      2155 => to_slv(opcode_type, 16#08#),
      2156 => to_slv(opcode_type, 16#05#),
      2157 => to_slv(opcode_type, 16#07#),
      2158 => to_slv(opcode_type, 16#0E#),
      2159 => to_slv(opcode_type, 16#0B#),
      2160 => to_slv(opcode_type, 16#06#),
      2161 => to_slv(opcode_type, 16#09#),
      2162 => to_slv(opcode_type, 16#0D#),
      2163 => to_slv(opcode_type, 16#0F#),
      2164 => to_slv(opcode_type, 16#09#),
      2165 => to_slv(opcode_type, 16#0D#),
      2166 => to_slv(opcode_type, 16#0E#),
      2167 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#09#),
      2177 => to_slv(opcode_type, 16#02#),
      2178 => to_slv(opcode_type, 16#07#),
      2179 => to_slv(opcode_type, 16#01#),
      2180 => to_slv(opcode_type, 16#0F#),
      2181 => to_slv(opcode_type, 16#09#),
      2182 => to_slv(opcode_type, 16#0F#),
      2183 => to_slv(opcode_type, 16#0D#),
      2184 => to_slv(opcode_type, 16#06#),
      2185 => to_slv(opcode_type, 16#08#),
      2186 => to_slv(opcode_type, 16#07#),
      2187 => to_slv(opcode_type, 16#0C#),
      2188 => to_slv(opcode_type, 16#0D#),
      2189 => to_slv(opcode_type, 16#08#),
      2190 => to_slv(opcode_type, 16#0B#),
      2191 => to_slv(opcode_type, 16#0F#),
      2192 => to_slv(opcode_type, 16#07#),
      2193 => to_slv(opcode_type, 16#09#),
      2194 => to_slv(opcode_type, 16#10#),
      2195 => to_slv(opcode_type, 16#0B#),
      2196 => to_slv(opcode_type, 16#09#),
      2197 => to_slv(opcode_type, 16#0B#),
      2198 => to_slv(opcode_type, 16#6E#),
      2199 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#06#),
      2209 => to_slv(opcode_type, 16#06#),
      2210 => to_slv(opcode_type, 16#06#),
      2211 => to_slv(opcode_type, 16#04#),
      2212 => to_slv(opcode_type, 16#0A#),
      2213 => to_slv(opcode_type, 16#04#),
      2214 => to_slv(opcode_type, 16#11#),
      2215 => to_slv(opcode_type, 16#03#),
      2216 => to_slv(opcode_type, 16#01#),
      2217 => to_slv(opcode_type, 16#11#),
      2218 => to_slv(opcode_type, 16#06#),
      2219 => to_slv(opcode_type, 16#09#),
      2220 => to_slv(opcode_type, 16#04#),
      2221 => to_slv(opcode_type, 16#0A#),
      2222 => to_slv(opcode_type, 16#03#),
      2223 => to_slv(opcode_type, 16#3C#),
      2224 => to_slv(opcode_type, 16#07#),
      2225 => to_slv(opcode_type, 16#06#),
      2226 => to_slv(opcode_type, 16#0B#),
      2227 => to_slv(opcode_type, 16#DA#),
      2228 => to_slv(opcode_type, 16#08#),
      2229 => to_slv(opcode_type, 16#11#),
      2230 => to_slv(opcode_type, 16#0B#),
      2231 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#02#),
      2242 => to_slv(opcode_type, 16#07#),
      2243 => to_slv(opcode_type, 16#08#),
      2244 => to_slv(opcode_type, 16#0F#),
      2245 => to_slv(opcode_type, 16#0A#),
      2246 => to_slv(opcode_type, 16#06#),
      2247 => to_slv(opcode_type, 16#0E#),
      2248 => to_slv(opcode_type, 16#0A#),
      2249 => to_slv(opcode_type, 16#09#),
      2250 => to_slv(opcode_type, 16#06#),
      2251 => to_slv(opcode_type, 16#04#),
      2252 => to_slv(opcode_type, 16#11#),
      2253 => to_slv(opcode_type, 16#06#),
      2254 => to_slv(opcode_type, 16#0F#),
      2255 => to_slv(opcode_type, 16#0F#),
      2256 => to_slv(opcode_type, 16#06#),
      2257 => to_slv(opcode_type, 16#07#),
      2258 => to_slv(opcode_type, 16#0E#),
      2259 => to_slv(opcode_type, 16#0E#),
      2260 => to_slv(opcode_type, 16#08#),
      2261 => to_slv(opcode_type, 16#74#),
      2262 => to_slv(opcode_type, 16#11#),
      2263 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#06#),
      2273 => to_slv(opcode_type, 16#01#),
      2274 => to_slv(opcode_type, 16#07#),
      2275 => to_slv(opcode_type, 16#05#),
      2276 => to_slv(opcode_type, 16#0C#),
      2277 => to_slv(opcode_type, 16#07#),
      2278 => to_slv(opcode_type, 16#10#),
      2279 => to_slv(opcode_type, 16#0B#),
      2280 => to_slv(opcode_type, 16#08#),
      2281 => to_slv(opcode_type, 16#08#),
      2282 => to_slv(opcode_type, 16#09#),
      2283 => to_slv(opcode_type, 16#0E#),
      2284 => to_slv(opcode_type, 16#10#),
      2285 => to_slv(opcode_type, 16#08#),
      2286 => to_slv(opcode_type, 16#4E#),
      2287 => to_slv(opcode_type, 16#0B#),
      2288 => to_slv(opcode_type, 16#08#),
      2289 => to_slv(opcode_type, 16#06#),
      2290 => to_slv(opcode_type, 16#0F#),
      2291 => to_slv(opcode_type, 16#10#),
      2292 => to_slv(opcode_type, 16#06#),
      2293 => to_slv(opcode_type, 16#C0#),
      2294 => to_slv(opcode_type, 16#0D#),
      2295 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#07#),
      2305 => to_slv(opcode_type, 16#07#),
      2306 => to_slv(opcode_type, 16#07#),
      2307 => to_slv(opcode_type, 16#03#),
      2308 => to_slv(opcode_type, 16#0B#),
      2309 => to_slv(opcode_type, 16#05#),
      2310 => to_slv(opcode_type, 16#0F#),
      2311 => to_slv(opcode_type, 16#04#),
      2312 => to_slv(opcode_type, 16#07#),
      2313 => to_slv(opcode_type, 16#10#),
      2314 => to_slv(opcode_type, 16#11#),
      2315 => to_slv(opcode_type, 16#08#),
      2316 => to_slv(opcode_type, 16#01#),
      2317 => to_slv(opcode_type, 16#09#),
      2318 => to_slv(opcode_type, 16#0F#),
      2319 => to_slv(opcode_type, 16#7F#),
      2320 => to_slv(opcode_type, 16#07#),
      2321 => to_slv(opcode_type, 16#06#),
      2322 => to_slv(opcode_type, 16#11#),
      2323 => to_slv(opcode_type, 16#0A#),
      2324 => to_slv(opcode_type, 16#09#),
      2325 => to_slv(opcode_type, 16#11#),
      2326 => to_slv(opcode_type, 16#0D#),
      2327 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#09#),
      2337 => to_slv(opcode_type, 16#03#),
      2338 => to_slv(opcode_type, 16#06#),
      2339 => to_slv(opcode_type, 16#01#),
      2340 => to_slv(opcode_type, 16#0A#),
      2341 => to_slv(opcode_type, 16#06#),
      2342 => to_slv(opcode_type, 16#0A#),
      2343 => to_slv(opcode_type, 16#0A#),
      2344 => to_slv(opcode_type, 16#08#),
      2345 => to_slv(opcode_type, 16#07#),
      2346 => to_slv(opcode_type, 16#08#),
      2347 => to_slv(opcode_type, 16#11#),
      2348 => to_slv(opcode_type, 16#11#),
      2349 => to_slv(opcode_type, 16#08#),
      2350 => to_slv(opcode_type, 16#0F#),
      2351 => to_slv(opcode_type, 16#10#),
      2352 => to_slv(opcode_type, 16#07#),
      2353 => to_slv(opcode_type, 16#07#),
      2354 => to_slv(opcode_type, 16#11#),
      2355 => to_slv(opcode_type, 16#0E#),
      2356 => to_slv(opcode_type, 16#07#),
      2357 => to_slv(opcode_type, 16#51#),
      2358 => to_slv(opcode_type, 16#0B#),
      2359 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#06#),
      2369 => to_slv(opcode_type, 16#09#),
      2370 => to_slv(opcode_type, 16#06#),
      2371 => to_slv(opcode_type, 16#04#),
      2372 => to_slv(opcode_type, 16#11#),
      2373 => to_slv(opcode_type, 16#07#),
      2374 => to_slv(opcode_type, 16#0F#),
      2375 => to_slv(opcode_type, 16#0F#),
      2376 => to_slv(opcode_type, 16#09#),
      2377 => to_slv(opcode_type, 16#08#),
      2378 => to_slv(opcode_type, 16#0A#),
      2379 => to_slv(opcode_type, 16#0F#),
      2380 => to_slv(opcode_type, 16#02#),
      2381 => to_slv(opcode_type, 16#0F#),
      2382 => to_slv(opcode_type, 16#07#),
      2383 => to_slv(opcode_type, 16#07#),
      2384 => to_slv(opcode_type, 16#04#),
      2385 => to_slv(opcode_type, 16#11#),
      2386 => to_slv(opcode_type, 16#04#),
      2387 => to_slv(opcode_type, 16#0A#),
      2388 => to_slv(opcode_type, 16#04#),
      2389 => to_slv(opcode_type, 16#03#),
      2390 => to_slv(opcode_type, 16#0F#),
      2391 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#09#),
      2401 => to_slv(opcode_type, 16#07#),
      2402 => to_slv(opcode_type, 16#04#),
      2403 => to_slv(opcode_type, 16#05#),
      2404 => to_slv(opcode_type, 16#0E#),
      2405 => to_slv(opcode_type, 16#03#),
      2406 => to_slv(opcode_type, 16#05#),
      2407 => to_slv(opcode_type, 16#0D#),
      2408 => to_slv(opcode_type, 16#08#),
      2409 => to_slv(opcode_type, 16#09#),
      2410 => to_slv(opcode_type, 16#09#),
      2411 => to_slv(opcode_type, 16#0C#),
      2412 => to_slv(opcode_type, 16#0E#),
      2413 => to_slv(opcode_type, 16#06#),
      2414 => to_slv(opcode_type, 16#0D#),
      2415 => to_slv(opcode_type, 16#0D#),
      2416 => to_slv(opcode_type, 16#08#),
      2417 => to_slv(opcode_type, 16#09#),
      2418 => to_slv(opcode_type, 16#0A#),
      2419 => to_slv(opcode_type, 16#0B#),
      2420 => to_slv(opcode_type, 16#07#),
      2421 => to_slv(opcode_type, 16#0C#),
      2422 => to_slv(opcode_type, 16#0A#),
      2423 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#07#),
      2433 => to_slv(opcode_type, 16#04#),
      2434 => to_slv(opcode_type, 16#08#),
      2435 => to_slv(opcode_type, 16#09#),
      2436 => to_slv(opcode_type, 16#0F#),
      2437 => to_slv(opcode_type, 16#0A#),
      2438 => to_slv(opcode_type, 16#06#),
      2439 => to_slv(opcode_type, 16#0A#),
      2440 => to_slv(opcode_type, 16#10#),
      2441 => to_slv(opcode_type, 16#07#),
      2442 => to_slv(opcode_type, 16#09#),
      2443 => to_slv(opcode_type, 16#08#),
      2444 => to_slv(opcode_type, 16#10#),
      2445 => to_slv(opcode_type, 16#11#),
      2446 => to_slv(opcode_type, 16#03#),
      2447 => to_slv(opcode_type, 16#0B#),
      2448 => to_slv(opcode_type, 16#08#),
      2449 => to_slv(opcode_type, 16#08#),
      2450 => to_slv(opcode_type, 16#0D#),
      2451 => to_slv(opcode_type, 16#0B#),
      2452 => to_slv(opcode_type, 16#06#),
      2453 => to_slv(opcode_type, 16#0B#),
      2454 => to_slv(opcode_type, 16#10#),
      2455 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#08#),
      2465 => to_slv(opcode_type, 16#07#),
      2466 => to_slv(opcode_type, 16#09#),
      2467 => to_slv(opcode_type, 16#03#),
      2468 => to_slv(opcode_type, 16#0A#),
      2469 => to_slv(opcode_type, 16#04#),
      2470 => to_slv(opcode_type, 16#C0#),
      2471 => to_slv(opcode_type, 16#02#),
      2472 => to_slv(opcode_type, 16#04#),
      2473 => to_slv(opcode_type, 16#CE#),
      2474 => to_slv(opcode_type, 16#06#),
      2475 => to_slv(opcode_type, 16#07#),
      2476 => to_slv(opcode_type, 16#02#),
      2477 => to_slv(opcode_type, 16#0D#),
      2478 => to_slv(opcode_type, 16#08#),
      2479 => to_slv(opcode_type, 16#0A#),
      2480 => to_slv(opcode_type, 16#11#),
      2481 => to_slv(opcode_type, 16#08#),
      2482 => to_slv(opcode_type, 16#06#),
      2483 => to_slv(opcode_type, 16#0F#),
      2484 => to_slv(opcode_type, 16#A7#),
      2485 => to_slv(opcode_type, 16#04#),
      2486 => to_slv(opcode_type, 16#0C#),
      2487 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#07#),
      2497 => to_slv(opcode_type, 16#09#),
      2498 => to_slv(opcode_type, 16#07#),
      2499 => to_slv(opcode_type, 16#09#),
      2500 => to_slv(opcode_type, 16#0E#),
      2501 => to_slv(opcode_type, 16#10#),
      2502 => to_slv(opcode_type, 16#04#),
      2503 => to_slv(opcode_type, 16#10#),
      2504 => to_slv(opcode_type, 16#05#),
      2505 => to_slv(opcode_type, 16#05#),
      2506 => to_slv(opcode_type, 16#0F#),
      2507 => to_slv(opcode_type, 16#07#),
      2508 => to_slv(opcode_type, 16#07#),
      2509 => to_slv(opcode_type, 16#03#),
      2510 => to_slv(opcode_type, 16#0C#),
      2511 => to_slv(opcode_type, 16#02#),
      2512 => to_slv(opcode_type, 16#0B#),
      2513 => to_slv(opcode_type, 16#09#),
      2514 => to_slv(opcode_type, 16#04#),
      2515 => to_slv(opcode_type, 16#0C#),
      2516 => to_slv(opcode_type, 16#07#),
      2517 => to_slv(opcode_type, 16#0E#),
      2518 => to_slv(opcode_type, 16#0C#),
      2519 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#04#),
      2530 => to_slv(opcode_type, 16#09#),
      2531 => to_slv(opcode_type, 16#05#),
      2532 => to_slv(opcode_type, 16#0B#),
      2533 => to_slv(opcode_type, 16#06#),
      2534 => to_slv(opcode_type, 16#0A#),
      2535 => to_slv(opcode_type, 16#0E#),
      2536 => to_slv(opcode_type, 16#07#),
      2537 => to_slv(opcode_type, 16#07#),
      2538 => to_slv(opcode_type, 16#08#),
      2539 => to_slv(opcode_type, 16#11#),
      2540 => to_slv(opcode_type, 16#0E#),
      2541 => to_slv(opcode_type, 16#08#),
      2542 => to_slv(opcode_type, 16#11#),
      2543 => to_slv(opcode_type, 16#0E#),
      2544 => to_slv(opcode_type, 16#09#),
      2545 => to_slv(opcode_type, 16#09#),
      2546 => to_slv(opcode_type, 16#14#),
      2547 => to_slv(opcode_type, 16#0D#),
      2548 => to_slv(opcode_type, 16#09#),
      2549 => to_slv(opcode_type, 16#F3#),
      2550 => to_slv(opcode_type, 16#0F#),
      2551 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#06#),
      2561 => to_slv(opcode_type, 16#02#),
      2562 => to_slv(opcode_type, 16#06#),
      2563 => to_slv(opcode_type, 16#06#),
      2564 => to_slv(opcode_type, 16#0F#),
      2565 => to_slv(opcode_type, 16#0B#),
      2566 => to_slv(opcode_type, 16#07#),
      2567 => to_slv(opcode_type, 16#0F#),
      2568 => to_slv(opcode_type, 16#0D#),
      2569 => to_slv(opcode_type, 16#06#),
      2570 => to_slv(opcode_type, 16#06#),
      2571 => to_slv(opcode_type, 16#02#),
      2572 => to_slv(opcode_type, 16#11#),
      2573 => to_slv(opcode_type, 16#06#),
      2574 => to_slv(opcode_type, 16#0E#),
      2575 => to_slv(opcode_type, 16#FB#),
      2576 => to_slv(opcode_type, 16#07#),
      2577 => to_slv(opcode_type, 16#09#),
      2578 => to_slv(opcode_type, 16#0B#),
      2579 => to_slv(opcode_type, 16#0E#),
      2580 => to_slv(opcode_type, 16#06#),
      2581 => to_slv(opcode_type, 16#0B#),
      2582 => to_slv(opcode_type, 16#DD#),
      2583 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#06#),
      2593 => to_slv(opcode_type, 16#04#),
      2594 => to_slv(opcode_type, 16#09#),
      2595 => to_slv(opcode_type, 16#06#),
      2596 => to_slv(opcode_type, 16#FB#),
      2597 => to_slv(opcode_type, 16#11#),
      2598 => to_slv(opcode_type, 16#08#),
      2599 => to_slv(opcode_type, 16#0D#),
      2600 => to_slv(opcode_type, 16#11#),
      2601 => to_slv(opcode_type, 16#09#),
      2602 => to_slv(opcode_type, 16#09#),
      2603 => to_slv(opcode_type, 16#04#),
      2604 => to_slv(opcode_type, 16#0A#),
      2605 => to_slv(opcode_type, 16#08#),
      2606 => to_slv(opcode_type, 16#0D#),
      2607 => to_slv(opcode_type, 16#11#),
      2608 => to_slv(opcode_type, 16#09#),
      2609 => to_slv(opcode_type, 16#08#),
      2610 => to_slv(opcode_type, 16#0E#),
      2611 => to_slv(opcode_type, 16#11#),
      2612 => to_slv(opcode_type, 16#07#),
      2613 => to_slv(opcode_type, 16#0F#),
      2614 => to_slv(opcode_type, 16#0B#),
      2615 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#06#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#01#),
      2627 => to_slv(opcode_type, 16#03#),
      2628 => to_slv(opcode_type, 16#6D#),
      2629 => to_slv(opcode_type, 16#08#),
      2630 => to_slv(opcode_type, 16#06#),
      2631 => to_slv(opcode_type, 16#0F#),
      2632 => to_slv(opcode_type, 16#0A#),
      2633 => to_slv(opcode_type, 16#02#),
      2634 => to_slv(opcode_type, 16#0D#),
      2635 => to_slv(opcode_type, 16#06#),
      2636 => to_slv(opcode_type, 16#01#),
      2637 => to_slv(opcode_type, 16#07#),
      2638 => to_slv(opcode_type, 16#0B#),
      2639 => to_slv(opcode_type, 16#0A#),
      2640 => to_slv(opcode_type, 16#09#),
      2641 => to_slv(opcode_type, 16#07#),
      2642 => to_slv(opcode_type, 16#0D#),
      2643 => to_slv(opcode_type, 16#10#),
      2644 => to_slv(opcode_type, 16#08#),
      2645 => to_slv(opcode_type, 16#71#),
      2646 => to_slv(opcode_type, 16#11#),
      2647 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#06#),
      2657 => to_slv(opcode_type, 16#08#),
      2658 => to_slv(opcode_type, 16#06#),
      2659 => to_slv(opcode_type, 16#02#),
      2660 => to_slv(opcode_type, 16#0F#),
      2661 => to_slv(opcode_type, 16#08#),
      2662 => to_slv(opcode_type, 16#0D#),
      2663 => to_slv(opcode_type, 16#0A#),
      2664 => to_slv(opcode_type, 16#02#),
      2665 => to_slv(opcode_type, 16#01#),
      2666 => to_slv(opcode_type, 16#0B#),
      2667 => to_slv(opcode_type, 16#08#),
      2668 => to_slv(opcode_type, 16#06#),
      2669 => to_slv(opcode_type, 16#01#),
      2670 => to_slv(opcode_type, 16#10#),
      2671 => to_slv(opcode_type, 16#03#),
      2672 => to_slv(opcode_type, 16#AD#),
      2673 => to_slv(opcode_type, 16#09#),
      2674 => to_slv(opcode_type, 16#05#),
      2675 => to_slv(opcode_type, 16#10#),
      2676 => to_slv(opcode_type, 16#07#),
      2677 => to_slv(opcode_type, 16#2E#),
      2678 => to_slv(opcode_type, 16#0A#),
      2679 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#09#),
      2689 => to_slv(opcode_type, 16#09#),
      2690 => to_slv(opcode_type, 16#03#),
      2691 => to_slv(opcode_type, 16#04#),
      2692 => to_slv(opcode_type, 16#0D#),
      2693 => to_slv(opcode_type, 16#05#),
      2694 => to_slv(opcode_type, 16#09#),
      2695 => to_slv(opcode_type, 16#10#),
      2696 => to_slv(opcode_type, 16#0C#),
      2697 => to_slv(opcode_type, 16#08#),
      2698 => to_slv(opcode_type, 16#09#),
      2699 => to_slv(opcode_type, 16#05#),
      2700 => to_slv(opcode_type, 16#0B#),
      2701 => to_slv(opcode_type, 16#09#),
      2702 => to_slv(opcode_type, 16#0A#),
      2703 => to_slv(opcode_type, 16#0B#),
      2704 => to_slv(opcode_type, 16#06#),
      2705 => to_slv(opcode_type, 16#06#),
      2706 => to_slv(opcode_type, 16#0B#),
      2707 => to_slv(opcode_type, 16#0D#),
      2708 => to_slv(opcode_type, 16#09#),
      2709 => to_slv(opcode_type, 16#0C#),
      2710 => to_slv(opcode_type, 16#0E#),
      2711 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#06#),
      2721 => to_slv(opcode_type, 16#01#),
      2722 => to_slv(opcode_type, 16#07#),
      2723 => to_slv(opcode_type, 16#08#),
      2724 => to_slv(opcode_type, 16#11#),
      2725 => to_slv(opcode_type, 16#0F#),
      2726 => to_slv(opcode_type, 16#02#),
      2727 => to_slv(opcode_type, 16#0E#),
      2728 => to_slv(opcode_type, 16#09#),
      2729 => to_slv(opcode_type, 16#09#),
      2730 => to_slv(opcode_type, 16#07#),
      2731 => to_slv(opcode_type, 16#10#),
      2732 => to_slv(opcode_type, 16#0D#),
      2733 => to_slv(opcode_type, 16#09#),
      2734 => to_slv(opcode_type, 16#0B#),
      2735 => to_slv(opcode_type, 16#0B#),
      2736 => to_slv(opcode_type, 16#07#),
      2737 => to_slv(opcode_type, 16#09#),
      2738 => to_slv(opcode_type, 16#10#),
      2739 => to_slv(opcode_type, 16#0C#),
      2740 => to_slv(opcode_type, 16#08#),
      2741 => to_slv(opcode_type, 16#0B#),
      2742 => to_slv(opcode_type, 16#0E#),
      2743 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#07#),
      2753 => to_slv(opcode_type, 16#04#),
      2754 => to_slv(opcode_type, 16#09#),
      2755 => to_slv(opcode_type, 16#03#),
      2756 => to_slv(opcode_type, 16#0D#),
      2757 => to_slv(opcode_type, 16#07#),
      2758 => to_slv(opcode_type, 16#11#),
      2759 => to_slv(opcode_type, 16#0B#),
      2760 => to_slv(opcode_type, 16#07#),
      2761 => to_slv(opcode_type, 16#08#),
      2762 => to_slv(opcode_type, 16#09#),
      2763 => to_slv(opcode_type, 16#11#),
      2764 => to_slv(opcode_type, 16#0F#),
      2765 => to_slv(opcode_type, 16#09#),
      2766 => to_slv(opcode_type, 16#0F#),
      2767 => to_slv(opcode_type, 16#11#),
      2768 => to_slv(opcode_type, 16#08#),
      2769 => to_slv(opcode_type, 16#07#),
      2770 => to_slv(opcode_type, 16#EA#),
      2771 => to_slv(opcode_type, 16#0D#),
      2772 => to_slv(opcode_type, 16#07#),
      2773 => to_slv(opcode_type, 16#0E#),
      2774 => to_slv(opcode_type, 16#0B#),
      2775 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#07#),
      2785 => to_slv(opcode_type, 16#08#),
      2786 => to_slv(opcode_type, 16#04#),
      2787 => to_slv(opcode_type, 16#09#),
      2788 => to_slv(opcode_type, 16#0D#),
      2789 => to_slv(opcode_type, 16#0E#),
      2790 => to_slv(opcode_type, 16#01#),
      2791 => to_slv(opcode_type, 16#03#),
      2792 => to_slv(opcode_type, 16#0C#),
      2793 => to_slv(opcode_type, 16#06#),
      2794 => to_slv(opcode_type, 16#07#),
      2795 => to_slv(opcode_type, 16#06#),
      2796 => to_slv(opcode_type, 16#0B#),
      2797 => to_slv(opcode_type, 16#11#),
      2798 => to_slv(opcode_type, 16#04#),
      2799 => to_slv(opcode_type, 16#0E#),
      2800 => to_slv(opcode_type, 16#07#),
      2801 => to_slv(opcode_type, 16#09#),
      2802 => to_slv(opcode_type, 16#0B#),
      2803 => to_slv(opcode_type, 16#11#),
      2804 => to_slv(opcode_type, 16#09#),
      2805 => to_slv(opcode_type, 16#0C#),
      2806 => to_slv(opcode_type, 16#0D#),
      2807 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#07#),
      2817 => to_slv(opcode_type, 16#01#),
      2818 => to_slv(opcode_type, 16#09#),
      2819 => to_slv(opcode_type, 16#07#),
      2820 => to_slv(opcode_type, 16#11#),
      2821 => to_slv(opcode_type, 16#11#),
      2822 => to_slv(opcode_type, 16#05#),
      2823 => to_slv(opcode_type, 16#0B#),
      2824 => to_slv(opcode_type, 16#09#),
      2825 => to_slv(opcode_type, 16#09#),
      2826 => to_slv(opcode_type, 16#09#),
      2827 => to_slv(opcode_type, 16#10#),
      2828 => to_slv(opcode_type, 16#0C#),
      2829 => to_slv(opcode_type, 16#08#),
      2830 => to_slv(opcode_type, 16#0B#),
      2831 => to_slv(opcode_type, 16#0E#),
      2832 => to_slv(opcode_type, 16#06#),
      2833 => to_slv(opcode_type, 16#07#),
      2834 => to_slv(opcode_type, 16#10#),
      2835 => to_slv(opcode_type, 16#0C#),
      2836 => to_slv(opcode_type, 16#09#),
      2837 => to_slv(opcode_type, 16#0B#),
      2838 => to_slv(opcode_type, 16#0B#),
      2839 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#09#),
      2849 => to_slv(opcode_type, 16#02#),
      2850 => to_slv(opcode_type, 16#06#),
      2851 => to_slv(opcode_type, 16#03#),
      2852 => to_slv(opcode_type, 16#0F#),
      2853 => to_slv(opcode_type, 16#09#),
      2854 => to_slv(opcode_type, 16#0E#),
      2855 => to_slv(opcode_type, 16#0B#),
      2856 => to_slv(opcode_type, 16#09#),
      2857 => to_slv(opcode_type, 16#06#),
      2858 => to_slv(opcode_type, 16#07#),
      2859 => to_slv(opcode_type, 16#10#),
      2860 => to_slv(opcode_type, 16#0B#),
      2861 => to_slv(opcode_type, 16#07#),
      2862 => to_slv(opcode_type, 16#0C#),
      2863 => to_slv(opcode_type, 16#0C#),
      2864 => to_slv(opcode_type, 16#08#),
      2865 => to_slv(opcode_type, 16#07#),
      2866 => to_slv(opcode_type, 16#0A#),
      2867 => to_slv(opcode_type, 16#0E#),
      2868 => to_slv(opcode_type, 16#06#),
      2869 => to_slv(opcode_type, 16#0E#),
      2870 => to_slv(opcode_type, 16#0F#),
      2871 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#07#),
      2881 => to_slv(opcode_type, 16#03#),
      2882 => to_slv(opcode_type, 16#06#),
      2883 => to_slv(opcode_type, 16#09#),
      2884 => to_slv(opcode_type, 16#10#),
      2885 => to_slv(opcode_type, 16#11#),
      2886 => to_slv(opcode_type, 16#03#),
      2887 => to_slv(opcode_type, 16#0C#),
      2888 => to_slv(opcode_type, 16#08#),
      2889 => to_slv(opcode_type, 16#08#),
      2890 => to_slv(opcode_type, 16#09#),
      2891 => to_slv(opcode_type, 16#0D#),
      2892 => to_slv(opcode_type, 16#C2#),
      2893 => to_slv(opcode_type, 16#06#),
      2894 => to_slv(opcode_type, 16#0C#),
      2895 => to_slv(opcode_type, 16#0D#),
      2896 => to_slv(opcode_type, 16#09#),
      2897 => to_slv(opcode_type, 16#06#),
      2898 => to_slv(opcode_type, 16#0F#),
      2899 => to_slv(opcode_type, 16#97#),
      2900 => to_slv(opcode_type, 16#06#),
      2901 => to_slv(opcode_type, 16#11#),
      2902 => to_slv(opcode_type, 16#0F#),
      2903 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#07#),
      2913 => to_slv(opcode_type, 16#05#),
      2914 => to_slv(opcode_type, 16#07#),
      2915 => to_slv(opcode_type, 16#09#),
      2916 => to_slv(opcode_type, 16#0C#),
      2917 => to_slv(opcode_type, 16#0D#),
      2918 => to_slv(opcode_type, 16#09#),
      2919 => to_slv(opcode_type, 16#0F#),
      2920 => to_slv(opcode_type, 16#ED#),
      2921 => to_slv(opcode_type, 16#06#),
      2922 => to_slv(opcode_type, 16#09#),
      2923 => to_slv(opcode_type, 16#03#),
      2924 => to_slv(opcode_type, 16#64#),
      2925 => to_slv(opcode_type, 16#07#),
      2926 => to_slv(opcode_type, 16#0F#),
      2927 => to_slv(opcode_type, 16#0F#),
      2928 => to_slv(opcode_type, 16#09#),
      2929 => to_slv(opcode_type, 16#08#),
      2930 => to_slv(opcode_type, 16#45#),
      2931 => to_slv(opcode_type, 16#0D#),
      2932 => to_slv(opcode_type, 16#07#),
      2933 => to_slv(opcode_type, 16#11#),
      2934 => to_slv(opcode_type, 16#0E#),
      2935 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#08#),
      2945 => to_slv(opcode_type, 16#01#),
      2946 => to_slv(opcode_type, 16#06#),
      2947 => to_slv(opcode_type, 16#03#),
      2948 => to_slv(opcode_type, 16#0F#),
      2949 => to_slv(opcode_type, 16#08#),
      2950 => to_slv(opcode_type, 16#0E#),
      2951 => to_slv(opcode_type, 16#0B#),
      2952 => to_slv(opcode_type, 16#07#),
      2953 => to_slv(opcode_type, 16#06#),
      2954 => to_slv(opcode_type, 16#07#),
      2955 => to_slv(opcode_type, 16#11#),
      2956 => to_slv(opcode_type, 16#0A#),
      2957 => to_slv(opcode_type, 16#07#),
      2958 => to_slv(opcode_type, 16#10#),
      2959 => to_slv(opcode_type, 16#11#),
      2960 => to_slv(opcode_type, 16#09#),
      2961 => to_slv(opcode_type, 16#08#),
      2962 => to_slv(opcode_type, 16#0A#),
      2963 => to_slv(opcode_type, 16#0F#),
      2964 => to_slv(opcode_type, 16#07#),
      2965 => to_slv(opcode_type, 16#0A#),
      2966 => to_slv(opcode_type, 16#0D#),
      2967 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#09#),
      2977 => to_slv(opcode_type, 16#07#),
      2978 => to_slv(opcode_type, 16#07#),
      2979 => to_slv(opcode_type, 16#03#),
      2980 => to_slv(opcode_type, 16#0A#),
      2981 => to_slv(opcode_type, 16#01#),
      2982 => to_slv(opcode_type, 16#0E#),
      2983 => to_slv(opcode_type, 16#03#),
      2984 => to_slv(opcode_type, 16#02#),
      2985 => to_slv(opcode_type, 16#11#),
      2986 => to_slv(opcode_type, 16#07#),
      2987 => to_slv(opcode_type, 16#07#),
      2988 => to_slv(opcode_type, 16#01#),
      2989 => to_slv(opcode_type, 16#0E#),
      2990 => to_slv(opcode_type, 16#02#),
      2991 => to_slv(opcode_type, 16#0B#),
      2992 => to_slv(opcode_type, 16#06#),
      2993 => to_slv(opcode_type, 16#09#),
      2994 => to_slv(opcode_type, 16#10#),
      2995 => to_slv(opcode_type, 16#FC#),
      2996 => to_slv(opcode_type, 16#07#),
      2997 => to_slv(opcode_type, 16#0A#),
      2998 => to_slv(opcode_type, 16#10#),
      2999 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#07#),
      3009 => to_slv(opcode_type, 16#06#),
      3010 => to_slv(opcode_type, 16#05#),
      3011 => to_slv(opcode_type, 16#04#),
      3012 => to_slv(opcode_type, 16#0C#),
      3013 => to_slv(opcode_type, 16#09#),
      3014 => to_slv(opcode_type, 16#08#),
      3015 => to_slv(opcode_type, 16#0E#),
      3016 => to_slv(opcode_type, 16#0B#),
      3017 => to_slv(opcode_type, 16#09#),
      3018 => to_slv(opcode_type, 16#0C#),
      3019 => to_slv(opcode_type, 16#11#),
      3020 => to_slv(opcode_type, 16#06#),
      3021 => to_slv(opcode_type, 16#04#),
      3022 => to_slv(opcode_type, 16#09#),
      3023 => to_slv(opcode_type, 16#11#),
      3024 => to_slv(opcode_type, 16#0B#),
      3025 => to_slv(opcode_type, 16#06#),
      3026 => to_slv(opcode_type, 16#04#),
      3027 => to_slv(opcode_type, 16#0D#),
      3028 => to_slv(opcode_type, 16#09#),
      3029 => to_slv(opcode_type, 16#0F#),
      3030 => to_slv(opcode_type, 16#10#),
      3031 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#09#),
      3041 => to_slv(opcode_type, 16#05#),
      3042 => to_slv(opcode_type, 16#06#),
      3043 => to_slv(opcode_type, 16#06#),
      3044 => to_slv(opcode_type, 16#0E#),
      3045 => to_slv(opcode_type, 16#11#),
      3046 => to_slv(opcode_type, 16#09#),
      3047 => to_slv(opcode_type, 16#0E#),
      3048 => to_slv(opcode_type, 16#0E#),
      3049 => to_slv(opcode_type, 16#07#),
      3050 => to_slv(opcode_type, 16#06#),
      3051 => to_slv(opcode_type, 16#05#),
      3052 => to_slv(opcode_type, 16#0B#),
      3053 => to_slv(opcode_type, 16#06#),
      3054 => to_slv(opcode_type, 16#0A#),
      3055 => to_slv(opcode_type, 16#0E#),
      3056 => to_slv(opcode_type, 16#09#),
      3057 => to_slv(opcode_type, 16#08#),
      3058 => to_slv(opcode_type, 16#0F#),
      3059 => to_slv(opcode_type, 16#0A#),
      3060 => to_slv(opcode_type, 16#06#),
      3061 => to_slv(opcode_type, 16#0A#),
      3062 => to_slv(opcode_type, 16#0E#),
      3063 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#06#),
      3073 => to_slv(opcode_type, 16#09#),
      3074 => to_slv(opcode_type, 16#09#),
      3075 => to_slv(opcode_type, 16#08#),
      3076 => to_slv(opcode_type, 16#0D#),
      3077 => to_slv(opcode_type, 16#0A#),
      3078 => to_slv(opcode_type, 16#02#),
      3079 => to_slv(opcode_type, 16#0E#),
      3080 => to_slv(opcode_type, 16#06#),
      3081 => to_slv(opcode_type, 16#06#),
      3082 => to_slv(opcode_type, 16#0B#),
      3083 => to_slv(opcode_type, 16#0F#),
      3084 => to_slv(opcode_type, 16#05#),
      3085 => to_slv(opcode_type, 16#11#),
      3086 => to_slv(opcode_type, 16#08#),
      3087 => to_slv(opcode_type, 16#01#),
      3088 => to_slv(opcode_type, 16#01#),
      3089 => to_slv(opcode_type, 16#0D#),
      3090 => to_slv(opcode_type, 16#07#),
      3091 => to_slv(opcode_type, 16#01#),
      3092 => to_slv(opcode_type, 16#0B#),
      3093 => to_slv(opcode_type, 16#03#),
      3094 => to_slv(opcode_type, 16#FA#),
      3095 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#09#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#08#),
      3107 => to_slv(opcode_type, 16#02#),
      3108 => to_slv(opcode_type, 16#0A#),
      3109 => to_slv(opcode_type, 16#03#),
      3110 => to_slv(opcode_type, 16#11#),
      3111 => to_slv(opcode_type, 16#06#),
      3112 => to_slv(opcode_type, 16#07#),
      3113 => to_slv(opcode_type, 16#10#),
      3114 => to_slv(opcode_type, 16#11#),
      3115 => to_slv(opcode_type, 16#02#),
      3116 => to_slv(opcode_type, 16#10#),
      3117 => to_slv(opcode_type, 16#07#),
      3118 => to_slv(opcode_type, 16#03#),
      3119 => to_slv(opcode_type, 16#05#),
      3120 => to_slv(opcode_type, 16#11#),
      3121 => to_slv(opcode_type, 16#07#),
      3122 => to_slv(opcode_type, 16#06#),
      3123 => to_slv(opcode_type, 16#0C#),
      3124 => to_slv(opcode_type, 16#0E#),
      3125 => to_slv(opcode_type, 16#04#),
      3126 => to_slv(opcode_type, 16#10#),
      3127 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#07#),
      3137 => to_slv(opcode_type, 16#03#),
      3138 => to_slv(opcode_type, 16#06#),
      3139 => to_slv(opcode_type, 16#01#),
      3140 => to_slv(opcode_type, 16#0C#),
      3141 => to_slv(opcode_type, 16#08#),
      3142 => to_slv(opcode_type, 16#0C#),
      3143 => to_slv(opcode_type, 16#11#),
      3144 => to_slv(opcode_type, 16#08#),
      3145 => to_slv(opcode_type, 16#06#),
      3146 => to_slv(opcode_type, 16#09#),
      3147 => to_slv(opcode_type, 16#0C#),
      3148 => to_slv(opcode_type, 16#18#),
      3149 => to_slv(opcode_type, 16#06#),
      3150 => to_slv(opcode_type, 16#11#),
      3151 => to_slv(opcode_type, 16#11#),
      3152 => to_slv(opcode_type, 16#07#),
      3153 => to_slv(opcode_type, 16#09#),
      3154 => to_slv(opcode_type, 16#0D#),
      3155 => to_slv(opcode_type, 16#11#),
      3156 => to_slv(opcode_type, 16#09#),
      3157 => to_slv(opcode_type, 16#BC#),
      3158 => to_slv(opcode_type, 16#11#),
      3159 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#06#),
      3169 => to_slv(opcode_type, 16#04#),
      3170 => to_slv(opcode_type, 16#09#),
      3171 => to_slv(opcode_type, 16#07#),
      3172 => to_slv(opcode_type, 16#0E#),
      3173 => to_slv(opcode_type, 16#10#),
      3174 => to_slv(opcode_type, 16#09#),
      3175 => to_slv(opcode_type, 16#0D#),
      3176 => to_slv(opcode_type, 16#0A#),
      3177 => to_slv(opcode_type, 16#08#),
      3178 => to_slv(opcode_type, 16#09#),
      3179 => to_slv(opcode_type, 16#05#),
      3180 => to_slv(opcode_type, 16#10#),
      3181 => to_slv(opcode_type, 16#06#),
      3182 => to_slv(opcode_type, 16#0E#),
      3183 => to_slv(opcode_type, 16#0C#),
      3184 => to_slv(opcode_type, 16#08#),
      3185 => to_slv(opcode_type, 16#07#),
      3186 => to_slv(opcode_type, 16#0E#),
      3187 => to_slv(opcode_type, 16#16#),
      3188 => to_slv(opcode_type, 16#09#),
      3189 => to_slv(opcode_type, 16#0D#),
      3190 => to_slv(opcode_type, 16#10#),
      3191 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#06#),
      3201 => to_slv(opcode_type, 16#08#),
      3202 => to_slv(opcode_type, 16#08#),
      3203 => to_slv(opcode_type, 16#02#),
      3204 => to_slv(opcode_type, 16#0F#),
      3205 => to_slv(opcode_type, 16#03#),
      3206 => to_slv(opcode_type, 16#0D#),
      3207 => to_slv(opcode_type, 16#01#),
      3208 => to_slv(opcode_type, 16#01#),
      3209 => to_slv(opcode_type, 16#0A#),
      3210 => to_slv(opcode_type, 16#09#),
      3211 => to_slv(opcode_type, 16#06#),
      3212 => to_slv(opcode_type, 16#08#),
      3213 => to_slv(opcode_type, 16#0D#),
      3214 => to_slv(opcode_type, 16#0B#),
      3215 => to_slv(opcode_type, 16#02#),
      3216 => to_slv(opcode_type, 16#0F#),
      3217 => to_slv(opcode_type, 16#06#),
      3218 => to_slv(opcode_type, 16#02#),
      3219 => to_slv(opcode_type, 16#11#),
      3220 => to_slv(opcode_type, 16#08#),
      3221 => to_slv(opcode_type, 16#0E#),
      3222 => to_slv(opcode_type, 16#0D#),
      3223 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#07#),
      3233 => to_slv(opcode_type, 16#02#),
      3234 => to_slv(opcode_type, 16#06#),
      3235 => to_slv(opcode_type, 16#05#),
      3236 => to_slv(opcode_type, 16#0E#),
      3237 => to_slv(opcode_type, 16#08#),
      3238 => to_slv(opcode_type, 16#10#),
      3239 => to_slv(opcode_type, 16#0F#),
      3240 => to_slv(opcode_type, 16#06#),
      3241 => to_slv(opcode_type, 16#09#),
      3242 => to_slv(opcode_type, 16#07#),
      3243 => to_slv(opcode_type, 16#0B#),
      3244 => to_slv(opcode_type, 16#0B#),
      3245 => to_slv(opcode_type, 16#08#),
      3246 => to_slv(opcode_type, 16#0E#),
      3247 => to_slv(opcode_type, 16#10#),
      3248 => to_slv(opcode_type, 16#09#),
      3249 => to_slv(opcode_type, 16#08#),
      3250 => to_slv(opcode_type, 16#0D#),
      3251 => to_slv(opcode_type, 16#29#),
      3252 => to_slv(opcode_type, 16#06#),
      3253 => to_slv(opcode_type, 16#0A#),
      3254 => to_slv(opcode_type, 16#0F#),
      3255 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#09#),
      3265 => to_slv(opcode_type, 16#01#),
      3266 => to_slv(opcode_type, 16#07#),
      3267 => to_slv(opcode_type, 16#01#),
      3268 => to_slv(opcode_type, 16#0C#),
      3269 => to_slv(opcode_type, 16#08#),
      3270 => to_slv(opcode_type, 16#0E#),
      3271 => to_slv(opcode_type, 16#0D#),
      3272 => to_slv(opcode_type, 16#09#),
      3273 => to_slv(opcode_type, 16#09#),
      3274 => to_slv(opcode_type, 16#08#),
      3275 => to_slv(opcode_type, 16#0A#),
      3276 => to_slv(opcode_type, 16#0E#),
      3277 => to_slv(opcode_type, 16#07#),
      3278 => to_slv(opcode_type, 16#11#),
      3279 => to_slv(opcode_type, 16#0B#),
      3280 => to_slv(opcode_type, 16#08#),
      3281 => to_slv(opcode_type, 16#09#),
      3282 => to_slv(opcode_type, 16#10#),
      3283 => to_slv(opcode_type, 16#0C#),
      3284 => to_slv(opcode_type, 16#08#),
      3285 => to_slv(opcode_type, 16#0A#),
      3286 => to_slv(opcode_type, 16#0A#),
      3287 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#09#),
      3297 => to_slv(opcode_type, 16#06#),
      3298 => to_slv(opcode_type, 16#07#),
      3299 => to_slv(opcode_type, 16#04#),
      3300 => to_slv(opcode_type, 16#0B#),
      3301 => to_slv(opcode_type, 16#06#),
      3302 => to_slv(opcode_type, 16#0B#),
      3303 => to_slv(opcode_type, 16#0D#),
      3304 => to_slv(opcode_type, 16#07#),
      3305 => to_slv(opcode_type, 16#02#),
      3306 => to_slv(opcode_type, 16#10#),
      3307 => to_slv(opcode_type, 16#04#),
      3308 => to_slv(opcode_type, 16#0F#),
      3309 => to_slv(opcode_type, 16#08#),
      3310 => to_slv(opcode_type, 16#05#),
      3311 => to_slv(opcode_type, 16#09#),
      3312 => to_slv(opcode_type, 16#0A#),
      3313 => to_slv(opcode_type, 16#10#),
      3314 => to_slv(opcode_type, 16#06#),
      3315 => to_slv(opcode_type, 16#06#),
      3316 => to_slv(opcode_type, 16#0F#),
      3317 => to_slv(opcode_type, 16#0C#),
      3318 => to_slv(opcode_type, 16#10#),
      3319 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#08#),
      3329 => to_slv(opcode_type, 16#08#),
      3330 => to_slv(opcode_type, 16#08#),
      3331 => to_slv(opcode_type, 16#01#),
      3332 => to_slv(opcode_type, 16#47#),
      3333 => to_slv(opcode_type, 16#08#),
      3334 => to_slv(opcode_type, 16#0A#),
      3335 => to_slv(opcode_type, 16#0E#),
      3336 => to_slv(opcode_type, 16#09#),
      3337 => to_slv(opcode_type, 16#01#),
      3338 => to_slv(opcode_type, 16#0B#),
      3339 => to_slv(opcode_type, 16#03#),
      3340 => to_slv(opcode_type, 16#0D#),
      3341 => to_slv(opcode_type, 16#08#),
      3342 => to_slv(opcode_type, 16#07#),
      3343 => to_slv(opcode_type, 16#01#),
      3344 => to_slv(opcode_type, 16#0B#),
      3345 => to_slv(opcode_type, 16#08#),
      3346 => to_slv(opcode_type, 16#11#),
      3347 => to_slv(opcode_type, 16#10#),
      3348 => to_slv(opcode_type, 16#07#),
      3349 => to_slv(opcode_type, 16#0C#),
      3350 => to_slv(opcode_type, 16#11#),
      3351 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#06#),
      3361 => to_slv(opcode_type, 16#06#),
      3362 => to_slv(opcode_type, 16#09#),
      3363 => to_slv(opcode_type, 16#02#),
      3364 => to_slv(opcode_type, 16#10#),
      3365 => to_slv(opcode_type, 16#05#),
      3366 => to_slv(opcode_type, 16#0A#),
      3367 => to_slv(opcode_type, 16#07#),
      3368 => to_slv(opcode_type, 16#02#),
      3369 => to_slv(opcode_type, 16#0A#),
      3370 => to_slv(opcode_type, 16#03#),
      3371 => to_slv(opcode_type, 16#0F#),
      3372 => to_slv(opcode_type, 16#09#),
      3373 => to_slv(opcode_type, 16#06#),
      3374 => to_slv(opcode_type, 16#07#),
      3375 => to_slv(opcode_type, 16#0E#),
      3376 => to_slv(opcode_type, 16#0F#),
      3377 => to_slv(opcode_type, 16#07#),
      3378 => to_slv(opcode_type, 16#0D#),
      3379 => to_slv(opcode_type, 16#0D#),
      3380 => to_slv(opcode_type, 16#01#),
      3381 => to_slv(opcode_type, 16#02#),
      3382 => to_slv(opcode_type, 16#0C#),
      3383 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#06#),
      3393 => to_slv(opcode_type, 16#07#),
      3394 => to_slv(opcode_type, 16#02#),
      3395 => to_slv(opcode_type, 16#06#),
      3396 => to_slv(opcode_type, 16#0E#),
      3397 => to_slv(opcode_type, 16#0F#),
      3398 => to_slv(opcode_type, 16#04#),
      3399 => to_slv(opcode_type, 16#06#),
      3400 => to_slv(opcode_type, 16#3D#),
      3401 => to_slv(opcode_type, 16#0E#),
      3402 => to_slv(opcode_type, 16#09#),
      3403 => to_slv(opcode_type, 16#07#),
      3404 => to_slv(opcode_type, 16#09#),
      3405 => to_slv(opcode_type, 16#0F#),
      3406 => to_slv(opcode_type, 16#11#),
      3407 => to_slv(opcode_type, 16#04#),
      3408 => to_slv(opcode_type, 16#0C#),
      3409 => to_slv(opcode_type, 16#09#),
      3410 => to_slv(opcode_type, 16#08#),
      3411 => to_slv(opcode_type, 16#0E#),
      3412 => to_slv(opcode_type, 16#0B#),
      3413 => to_slv(opcode_type, 16#04#),
      3414 => to_slv(opcode_type, 16#0A#),
      3415 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#06#),
      3425 => to_slv(opcode_type, 16#08#),
      3426 => to_slv(opcode_type, 16#05#),
      3427 => to_slv(opcode_type, 16#04#),
      3428 => to_slv(opcode_type, 16#0E#),
      3429 => to_slv(opcode_type, 16#03#),
      3430 => to_slv(opcode_type, 16#03#),
      3431 => to_slv(opcode_type, 16#32#),
      3432 => to_slv(opcode_type, 16#06#),
      3433 => to_slv(opcode_type, 16#09#),
      3434 => to_slv(opcode_type, 16#06#),
      3435 => to_slv(opcode_type, 16#0A#),
      3436 => to_slv(opcode_type, 16#0C#),
      3437 => to_slv(opcode_type, 16#09#),
      3438 => to_slv(opcode_type, 16#10#),
      3439 => to_slv(opcode_type, 16#86#),
      3440 => to_slv(opcode_type, 16#07#),
      3441 => to_slv(opcode_type, 16#06#),
      3442 => to_slv(opcode_type, 16#44#),
      3443 => to_slv(opcode_type, 16#0D#),
      3444 => to_slv(opcode_type, 16#07#),
      3445 => to_slv(opcode_type, 16#0A#),
      3446 => to_slv(opcode_type, 16#0E#),
      3447 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#09#),
      3457 => to_slv(opcode_type, 16#03#),
      3458 => to_slv(opcode_type, 16#07#),
      3459 => to_slv(opcode_type, 16#04#),
      3460 => to_slv(opcode_type, 16#10#),
      3461 => to_slv(opcode_type, 16#07#),
      3462 => to_slv(opcode_type, 16#0E#),
      3463 => to_slv(opcode_type, 16#0C#),
      3464 => to_slv(opcode_type, 16#07#),
      3465 => to_slv(opcode_type, 16#09#),
      3466 => to_slv(opcode_type, 16#06#),
      3467 => to_slv(opcode_type, 16#0E#),
      3468 => to_slv(opcode_type, 16#0E#),
      3469 => to_slv(opcode_type, 16#08#),
      3470 => to_slv(opcode_type, 16#0A#),
      3471 => to_slv(opcode_type, 16#0B#),
      3472 => to_slv(opcode_type, 16#07#),
      3473 => to_slv(opcode_type, 16#08#),
      3474 => to_slv(opcode_type, 16#10#),
      3475 => to_slv(opcode_type, 16#0E#),
      3476 => to_slv(opcode_type, 16#09#),
      3477 => to_slv(opcode_type, 16#0C#),
      3478 => to_slv(opcode_type, 16#0E#),
      3479 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#09#),
      3489 => to_slv(opcode_type, 16#08#),
      3490 => to_slv(opcode_type, 16#07#),
      3491 => to_slv(opcode_type, 16#05#),
      3492 => to_slv(opcode_type, 16#10#),
      3493 => to_slv(opcode_type, 16#01#),
      3494 => to_slv(opcode_type, 16#10#),
      3495 => to_slv(opcode_type, 16#01#),
      3496 => to_slv(opcode_type, 16#07#),
      3497 => to_slv(opcode_type, 16#11#),
      3498 => to_slv(opcode_type, 16#0C#),
      3499 => to_slv(opcode_type, 16#08#),
      3500 => to_slv(opcode_type, 16#09#),
      3501 => to_slv(opcode_type, 16#08#),
      3502 => to_slv(opcode_type, 16#0B#),
      3503 => to_slv(opcode_type, 16#0F#),
      3504 => to_slv(opcode_type, 16#01#),
      3505 => to_slv(opcode_type, 16#3D#),
      3506 => to_slv(opcode_type, 16#08#),
      3507 => to_slv(opcode_type, 16#07#),
      3508 => to_slv(opcode_type, 16#10#),
      3509 => to_slv(opcode_type, 16#0C#),
      3510 => to_slv(opcode_type, 16#0A#),
      3511 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#07#),
      3521 => to_slv(opcode_type, 16#02#),
      3522 => to_slv(opcode_type, 16#07#),
      3523 => to_slv(opcode_type, 16#08#),
      3524 => to_slv(opcode_type, 16#0B#),
      3525 => to_slv(opcode_type, 16#11#),
      3526 => to_slv(opcode_type, 16#02#),
      3527 => to_slv(opcode_type, 16#0F#),
      3528 => to_slv(opcode_type, 16#08#),
      3529 => to_slv(opcode_type, 16#06#),
      3530 => to_slv(opcode_type, 16#07#),
      3531 => to_slv(opcode_type, 16#63#),
      3532 => to_slv(opcode_type, 16#0C#),
      3533 => to_slv(opcode_type, 16#08#),
      3534 => to_slv(opcode_type, 16#0A#),
      3535 => to_slv(opcode_type, 16#10#),
      3536 => to_slv(opcode_type, 16#08#),
      3537 => to_slv(opcode_type, 16#06#),
      3538 => to_slv(opcode_type, 16#0A#),
      3539 => to_slv(opcode_type, 16#0F#),
      3540 => to_slv(opcode_type, 16#09#),
      3541 => to_slv(opcode_type, 16#0A#),
      3542 => to_slv(opcode_type, 16#0A#),
      3543 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#06#),
      3553 => to_slv(opcode_type, 16#06#),
      3554 => to_slv(opcode_type, 16#01#),
      3555 => to_slv(opcode_type, 16#08#),
      3556 => to_slv(opcode_type, 16#0F#),
      3557 => to_slv(opcode_type, 16#FF#),
      3558 => to_slv(opcode_type, 16#01#),
      3559 => to_slv(opcode_type, 16#05#),
      3560 => to_slv(opcode_type, 16#0C#),
      3561 => to_slv(opcode_type, 16#06#),
      3562 => to_slv(opcode_type, 16#07#),
      3563 => to_slv(opcode_type, 16#04#),
      3564 => to_slv(opcode_type, 16#0D#),
      3565 => to_slv(opcode_type, 16#07#),
      3566 => to_slv(opcode_type, 16#10#),
      3567 => to_slv(opcode_type, 16#10#),
      3568 => to_slv(opcode_type, 16#06#),
      3569 => to_slv(opcode_type, 16#07#),
      3570 => to_slv(opcode_type, 16#0B#),
      3571 => to_slv(opcode_type, 16#0A#),
      3572 => to_slv(opcode_type, 16#09#),
      3573 => to_slv(opcode_type, 16#0C#),
      3574 => to_slv(opcode_type, 16#0B#),
      3575 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#09#),
      3585 => to_slv(opcode_type, 16#06#),
      3586 => to_slv(opcode_type, 16#06#),
      3587 => to_slv(opcode_type, 16#08#),
      3588 => to_slv(opcode_type, 16#11#),
      3589 => to_slv(opcode_type, 16#0D#),
      3590 => to_slv(opcode_type, 16#02#),
      3591 => to_slv(opcode_type, 16#10#),
      3592 => to_slv(opcode_type, 16#07#),
      3593 => to_slv(opcode_type, 16#02#),
      3594 => to_slv(opcode_type, 16#0A#),
      3595 => to_slv(opcode_type, 16#03#),
      3596 => to_slv(opcode_type, 16#0D#),
      3597 => to_slv(opcode_type, 16#08#),
      3598 => to_slv(opcode_type, 16#05#),
      3599 => to_slv(opcode_type, 16#07#),
      3600 => to_slv(opcode_type, 16#0B#),
      3601 => to_slv(opcode_type, 16#11#),
      3602 => to_slv(opcode_type, 16#06#),
      3603 => to_slv(opcode_type, 16#03#),
      3604 => to_slv(opcode_type, 16#0F#),
      3605 => to_slv(opcode_type, 16#05#),
      3606 => to_slv(opcode_type, 16#0F#),
      3607 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#07#),
      3617 => to_slv(opcode_type, 16#02#),
      3618 => to_slv(opcode_type, 16#08#),
      3619 => to_slv(opcode_type, 16#07#),
      3620 => to_slv(opcode_type, 16#11#),
      3621 => to_slv(opcode_type, 16#11#),
      3622 => to_slv(opcode_type, 16#08#),
      3623 => to_slv(opcode_type, 16#CA#),
      3624 => to_slv(opcode_type, 16#0A#),
      3625 => to_slv(opcode_type, 16#07#),
      3626 => to_slv(opcode_type, 16#06#),
      3627 => to_slv(opcode_type, 16#01#),
      3628 => to_slv(opcode_type, 16#0C#),
      3629 => to_slv(opcode_type, 16#07#),
      3630 => to_slv(opcode_type, 16#0C#),
      3631 => to_slv(opcode_type, 16#0C#),
      3632 => to_slv(opcode_type, 16#08#),
      3633 => to_slv(opcode_type, 16#08#),
      3634 => to_slv(opcode_type, 16#0A#),
      3635 => to_slv(opcode_type, 16#0C#),
      3636 => to_slv(opcode_type, 16#06#),
      3637 => to_slv(opcode_type, 16#0B#),
      3638 => to_slv(opcode_type, 16#0F#),
      3639 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#07#),
      3649 => to_slv(opcode_type, 16#01#),
      3650 => to_slv(opcode_type, 16#07#),
      3651 => to_slv(opcode_type, 16#09#),
      3652 => to_slv(opcode_type, 16#0D#),
      3653 => to_slv(opcode_type, 16#10#),
      3654 => to_slv(opcode_type, 16#09#),
      3655 => to_slv(opcode_type, 16#0D#),
      3656 => to_slv(opcode_type, 16#0A#),
      3657 => to_slv(opcode_type, 16#08#),
      3658 => to_slv(opcode_type, 16#09#),
      3659 => to_slv(opcode_type, 16#07#),
      3660 => to_slv(opcode_type, 16#0F#),
      3661 => to_slv(opcode_type, 16#0A#),
      3662 => to_slv(opcode_type, 16#08#),
      3663 => to_slv(opcode_type, 16#0D#),
      3664 => to_slv(opcode_type, 16#EF#),
      3665 => to_slv(opcode_type, 16#06#),
      3666 => to_slv(opcode_type, 16#02#),
      3667 => to_slv(opcode_type, 16#0B#),
      3668 => to_slv(opcode_type, 16#07#),
      3669 => to_slv(opcode_type, 16#0F#),
      3670 => to_slv(opcode_type, 16#39#),
      3671 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#09#),
      3681 => to_slv(opcode_type, 16#04#),
      3682 => to_slv(opcode_type, 16#07#),
      3683 => to_slv(opcode_type, 16#05#),
      3684 => to_slv(opcode_type, 16#0B#),
      3685 => to_slv(opcode_type, 16#06#),
      3686 => to_slv(opcode_type, 16#0B#),
      3687 => to_slv(opcode_type, 16#0F#),
      3688 => to_slv(opcode_type, 16#06#),
      3689 => to_slv(opcode_type, 16#09#),
      3690 => to_slv(opcode_type, 16#09#),
      3691 => to_slv(opcode_type, 16#10#),
      3692 => to_slv(opcode_type, 16#0D#),
      3693 => to_slv(opcode_type, 16#06#),
      3694 => to_slv(opcode_type, 16#11#),
      3695 => to_slv(opcode_type, 16#0F#),
      3696 => to_slv(opcode_type, 16#07#),
      3697 => to_slv(opcode_type, 16#08#),
      3698 => to_slv(opcode_type, 16#10#),
      3699 => to_slv(opcode_type, 16#10#),
      3700 => to_slv(opcode_type, 16#09#),
      3701 => to_slv(opcode_type, 16#0F#),
      3702 => to_slv(opcode_type, 16#11#),
      3703 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#07#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#04#),
      3715 => to_slv(opcode_type, 16#04#),
      3716 => to_slv(opcode_type, 16#10#),
      3717 => to_slv(opcode_type, 16#01#),
      3718 => to_slv(opcode_type, 16#04#),
      3719 => to_slv(opcode_type, 16#10#),
      3720 => to_slv(opcode_type, 16#07#),
      3721 => to_slv(opcode_type, 16#09#),
      3722 => to_slv(opcode_type, 16#07#),
      3723 => to_slv(opcode_type, 16#0C#),
      3724 => to_slv(opcode_type, 16#10#),
      3725 => to_slv(opcode_type, 16#06#),
      3726 => to_slv(opcode_type, 16#0D#),
      3727 => to_slv(opcode_type, 16#0A#),
      3728 => to_slv(opcode_type, 16#08#),
      3729 => to_slv(opcode_type, 16#06#),
      3730 => to_slv(opcode_type, 16#0D#),
      3731 => to_slv(opcode_type, 16#11#),
      3732 => to_slv(opcode_type, 16#08#),
      3733 => to_slv(opcode_type, 16#11#),
      3734 => to_slv(opcode_type, 16#0E#),
      3735 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#08#),
      3745 => to_slv(opcode_type, 16#06#),
      3746 => to_slv(opcode_type, 16#05#),
      3747 => to_slv(opcode_type, 16#08#),
      3748 => to_slv(opcode_type, 16#0B#),
      3749 => to_slv(opcode_type, 16#0B#),
      3750 => to_slv(opcode_type, 16#01#),
      3751 => to_slv(opcode_type, 16#08#),
      3752 => to_slv(opcode_type, 16#11#),
      3753 => to_slv(opcode_type, 16#0E#),
      3754 => to_slv(opcode_type, 16#07#),
      3755 => to_slv(opcode_type, 16#07#),
      3756 => to_slv(opcode_type, 16#08#),
      3757 => to_slv(opcode_type, 16#0D#),
      3758 => to_slv(opcode_type, 16#7D#),
      3759 => to_slv(opcode_type, 16#02#),
      3760 => to_slv(opcode_type, 16#0F#),
      3761 => to_slv(opcode_type, 16#09#),
      3762 => to_slv(opcode_type, 16#05#),
      3763 => to_slv(opcode_type, 16#0D#),
      3764 => to_slv(opcode_type, 16#09#),
      3765 => to_slv(opcode_type, 16#0F#),
      3766 => to_slv(opcode_type, 16#0C#),
      3767 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#09#),
      3777 => to_slv(opcode_type, 16#06#),
      3778 => to_slv(opcode_type, 16#07#),
      3779 => to_slv(opcode_type, 16#06#),
      3780 => to_slv(opcode_type, 16#10#),
      3781 => to_slv(opcode_type, 16#0A#),
      3782 => to_slv(opcode_type, 16#04#),
      3783 => to_slv(opcode_type, 16#0E#),
      3784 => to_slv(opcode_type, 16#05#),
      3785 => to_slv(opcode_type, 16#02#),
      3786 => to_slv(opcode_type, 16#0B#),
      3787 => to_slv(opcode_type, 16#09#),
      3788 => to_slv(opcode_type, 16#06#),
      3789 => to_slv(opcode_type, 16#09#),
      3790 => to_slv(opcode_type, 16#0C#),
      3791 => to_slv(opcode_type, 16#F1#),
      3792 => to_slv(opcode_type, 16#03#),
      3793 => to_slv(opcode_type, 16#0C#),
      3794 => to_slv(opcode_type, 16#09#),
      3795 => to_slv(opcode_type, 16#07#),
      3796 => to_slv(opcode_type, 16#0F#),
      3797 => to_slv(opcode_type, 16#10#),
      3798 => to_slv(opcode_type, 16#0D#),
      3799 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#06#),
      3809 => to_slv(opcode_type, 16#06#),
      3810 => to_slv(opcode_type, 16#09#),
      3811 => to_slv(opcode_type, 16#06#),
      3812 => to_slv(opcode_type, 16#F5#),
      3813 => to_slv(opcode_type, 16#11#),
      3814 => to_slv(opcode_type, 16#01#),
      3815 => to_slv(opcode_type, 16#0D#),
      3816 => to_slv(opcode_type, 16#05#),
      3817 => to_slv(opcode_type, 16#03#),
      3818 => to_slv(opcode_type, 16#10#),
      3819 => to_slv(opcode_type, 16#09#),
      3820 => to_slv(opcode_type, 16#03#),
      3821 => to_slv(opcode_type, 16#08#),
      3822 => to_slv(opcode_type, 16#0F#),
      3823 => to_slv(opcode_type, 16#11#),
      3824 => to_slv(opcode_type, 16#09#),
      3825 => to_slv(opcode_type, 16#06#),
      3826 => to_slv(opcode_type, 16#0A#),
      3827 => to_slv(opcode_type, 16#11#),
      3828 => to_slv(opcode_type, 16#08#),
      3829 => to_slv(opcode_type, 16#0F#),
      3830 => to_slv(opcode_type, 16#0C#),
      3831 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#06#),
      3841 => to_slv(opcode_type, 16#05#),
      3842 => to_slv(opcode_type, 16#09#),
      3843 => to_slv(opcode_type, 16#02#),
      3844 => to_slv(opcode_type, 16#11#),
      3845 => to_slv(opcode_type, 16#08#),
      3846 => to_slv(opcode_type, 16#0A#),
      3847 => to_slv(opcode_type, 16#34#),
      3848 => to_slv(opcode_type, 16#07#),
      3849 => to_slv(opcode_type, 16#08#),
      3850 => to_slv(opcode_type, 16#08#),
      3851 => to_slv(opcode_type, 16#0A#),
      3852 => to_slv(opcode_type, 16#0E#),
      3853 => to_slv(opcode_type, 16#07#),
      3854 => to_slv(opcode_type, 16#0B#),
      3855 => to_slv(opcode_type, 16#0D#),
      3856 => to_slv(opcode_type, 16#06#),
      3857 => to_slv(opcode_type, 16#07#),
      3858 => to_slv(opcode_type, 16#0B#),
      3859 => to_slv(opcode_type, 16#0B#),
      3860 => to_slv(opcode_type, 16#08#),
      3861 => to_slv(opcode_type, 16#0B#),
      3862 => to_slv(opcode_type, 16#0A#),
      3863 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#09#),
      3873 => to_slv(opcode_type, 16#08#),
      3874 => to_slv(opcode_type, 16#02#),
      3875 => to_slv(opcode_type, 16#08#),
      3876 => to_slv(opcode_type, 16#0F#),
      3877 => to_slv(opcode_type, 16#8B#),
      3878 => to_slv(opcode_type, 16#03#),
      3879 => to_slv(opcode_type, 16#06#),
      3880 => to_slv(opcode_type, 16#0F#),
      3881 => to_slv(opcode_type, 16#0D#),
      3882 => to_slv(opcode_type, 16#09#),
      3883 => to_slv(opcode_type, 16#07#),
      3884 => to_slv(opcode_type, 16#01#),
      3885 => to_slv(opcode_type, 16#0B#),
      3886 => to_slv(opcode_type, 16#07#),
      3887 => to_slv(opcode_type, 16#0D#),
      3888 => to_slv(opcode_type, 16#0D#),
      3889 => to_slv(opcode_type, 16#08#),
      3890 => to_slv(opcode_type, 16#04#),
      3891 => to_slv(opcode_type, 16#11#),
      3892 => to_slv(opcode_type, 16#06#),
      3893 => to_slv(opcode_type, 16#10#),
      3894 => to_slv(opcode_type, 16#0C#),
      3895 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#08#),
      3905 => to_slv(opcode_type, 16#01#),
      3906 => to_slv(opcode_type, 16#07#),
      3907 => to_slv(opcode_type, 16#07#),
      3908 => to_slv(opcode_type, 16#0A#),
      3909 => to_slv(opcode_type, 16#0F#),
      3910 => to_slv(opcode_type, 16#02#),
      3911 => to_slv(opcode_type, 16#11#),
      3912 => to_slv(opcode_type, 16#07#),
      3913 => to_slv(opcode_type, 16#06#),
      3914 => to_slv(opcode_type, 16#09#),
      3915 => to_slv(opcode_type, 16#0D#),
      3916 => to_slv(opcode_type, 16#0A#),
      3917 => to_slv(opcode_type, 16#07#),
      3918 => to_slv(opcode_type, 16#B9#),
      3919 => to_slv(opcode_type, 16#11#),
      3920 => to_slv(opcode_type, 16#08#),
      3921 => to_slv(opcode_type, 16#09#),
      3922 => to_slv(opcode_type, 16#0C#),
      3923 => to_slv(opcode_type, 16#0E#),
      3924 => to_slv(opcode_type, 16#06#),
      3925 => to_slv(opcode_type, 16#11#),
      3926 => to_slv(opcode_type, 16#0A#),
      3927 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#08#),
      3937 => to_slv(opcode_type, 16#01#),
      3938 => to_slv(opcode_type, 16#09#),
      3939 => to_slv(opcode_type, 16#03#),
      3940 => to_slv(opcode_type, 16#0B#),
      3941 => to_slv(opcode_type, 16#09#),
      3942 => to_slv(opcode_type, 16#0A#),
      3943 => to_slv(opcode_type, 16#0B#),
      3944 => to_slv(opcode_type, 16#08#),
      3945 => to_slv(opcode_type, 16#06#),
      3946 => to_slv(opcode_type, 16#09#),
      3947 => to_slv(opcode_type, 16#0C#),
      3948 => to_slv(opcode_type, 16#0D#),
      3949 => to_slv(opcode_type, 16#07#),
      3950 => to_slv(opcode_type, 16#0F#),
      3951 => to_slv(opcode_type, 16#0E#),
      3952 => to_slv(opcode_type, 16#07#),
      3953 => to_slv(opcode_type, 16#07#),
      3954 => to_slv(opcode_type, 16#0C#),
      3955 => to_slv(opcode_type, 16#10#),
      3956 => to_slv(opcode_type, 16#06#),
      3957 => to_slv(opcode_type, 16#11#),
      3958 => to_slv(opcode_type, 16#5E#),
      3959 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#08#),
      3969 => to_slv(opcode_type, 16#01#),
      3970 => to_slv(opcode_type, 16#08#),
      3971 => to_slv(opcode_type, 16#08#),
      3972 => to_slv(opcode_type, 16#0E#),
      3973 => to_slv(opcode_type, 16#46#),
      3974 => to_slv(opcode_type, 16#04#),
      3975 => to_slv(opcode_type, 16#0C#),
      3976 => to_slv(opcode_type, 16#06#),
      3977 => to_slv(opcode_type, 16#08#),
      3978 => to_slv(opcode_type, 16#09#),
      3979 => to_slv(opcode_type, 16#10#),
      3980 => to_slv(opcode_type, 16#0A#),
      3981 => to_slv(opcode_type, 16#09#),
      3982 => to_slv(opcode_type, 16#0A#),
      3983 => to_slv(opcode_type, 16#0F#),
      3984 => to_slv(opcode_type, 16#08#),
      3985 => to_slv(opcode_type, 16#07#),
      3986 => to_slv(opcode_type, 16#0C#),
      3987 => to_slv(opcode_type, 16#0A#),
      3988 => to_slv(opcode_type, 16#08#),
      3989 => to_slv(opcode_type, 16#0C#),
      3990 => to_slv(opcode_type, 16#0B#),
      3991 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#06#),
      4001 => to_slv(opcode_type, 16#09#),
      4002 => to_slv(opcode_type, 16#02#),
      4003 => to_slv(opcode_type, 16#06#),
      4004 => to_slv(opcode_type, 16#0F#),
      4005 => to_slv(opcode_type, 16#0D#),
      4006 => to_slv(opcode_type, 16#07#),
      4007 => to_slv(opcode_type, 16#07#),
      4008 => to_slv(opcode_type, 16#0B#),
      4009 => to_slv(opcode_type, 16#0A#),
      4010 => to_slv(opcode_type, 16#06#),
      4011 => to_slv(opcode_type, 16#83#),
      4012 => to_slv(opcode_type, 16#0C#),
      4013 => to_slv(opcode_type, 16#08#),
      4014 => to_slv(opcode_type, 16#09#),
      4015 => to_slv(opcode_type, 16#01#),
      4016 => to_slv(opcode_type, 16#0D#),
      4017 => to_slv(opcode_type, 16#09#),
      4018 => to_slv(opcode_type, 16#0C#),
      4019 => to_slv(opcode_type, 16#0F#),
      4020 => to_slv(opcode_type, 16#02#),
      4021 => to_slv(opcode_type, 16#05#),
      4022 => to_slv(opcode_type, 16#0E#),
      4023 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#07#),
      4033 => to_slv(opcode_type, 16#02#),
      4034 => to_slv(opcode_type, 16#09#),
      4035 => to_slv(opcode_type, 16#05#),
      4036 => to_slv(opcode_type, 16#0D#),
      4037 => to_slv(opcode_type, 16#09#),
      4038 => to_slv(opcode_type, 16#0D#),
      4039 => to_slv(opcode_type, 16#0C#),
      4040 => to_slv(opcode_type, 16#06#),
      4041 => to_slv(opcode_type, 16#08#),
      4042 => to_slv(opcode_type, 16#09#),
      4043 => to_slv(opcode_type, 16#0B#),
      4044 => to_slv(opcode_type, 16#0B#),
      4045 => to_slv(opcode_type, 16#08#),
      4046 => to_slv(opcode_type, 16#0F#),
      4047 => to_slv(opcode_type, 16#0F#),
      4048 => to_slv(opcode_type, 16#09#),
      4049 => to_slv(opcode_type, 16#08#),
      4050 => to_slv(opcode_type, 16#0C#),
      4051 => to_slv(opcode_type, 16#CB#),
      4052 => to_slv(opcode_type, 16#07#),
      4053 => to_slv(opcode_type, 16#0E#),
      4054 => to_slv(opcode_type, 16#10#),
      4055 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#08#),
      4065 => to_slv(opcode_type, 16#05#),
      4066 => to_slv(opcode_type, 16#08#),
      4067 => to_slv(opcode_type, 16#03#),
      4068 => to_slv(opcode_type, 16#0C#),
      4069 => to_slv(opcode_type, 16#06#),
      4070 => to_slv(opcode_type, 16#0A#),
      4071 => to_slv(opcode_type, 16#0C#),
      4072 => to_slv(opcode_type, 16#09#),
      4073 => to_slv(opcode_type, 16#08#),
      4074 => to_slv(opcode_type, 16#06#),
      4075 => to_slv(opcode_type, 16#11#),
      4076 => to_slv(opcode_type, 16#11#),
      4077 => to_slv(opcode_type, 16#06#),
      4078 => to_slv(opcode_type, 16#11#),
      4079 => to_slv(opcode_type, 16#0B#),
      4080 => to_slv(opcode_type, 16#09#),
      4081 => to_slv(opcode_type, 16#06#),
      4082 => to_slv(opcode_type, 16#10#),
      4083 => to_slv(opcode_type, 16#0D#),
      4084 => to_slv(opcode_type, 16#08#),
      4085 => to_slv(opcode_type, 16#0C#),
      4086 => to_slv(opcode_type, 16#11#),
      4087 to 4095 => (others => '0')
  ),

    -- Bin `24`...
    23 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#07#),
      1 => to_slv(opcode_type, 16#04#),
      2 => to_slv(opcode_type, 16#09#),
      3 => to_slv(opcode_type, 16#08#),
      4 => to_slv(opcode_type, 16#81#),
      5 => to_slv(opcode_type, 16#0E#),
      6 => to_slv(opcode_type, 16#08#),
      7 => to_slv(opcode_type, 16#0F#),
      8 => to_slv(opcode_type, 16#11#),
      9 => to_slv(opcode_type, 16#08#),
      10 => to_slv(opcode_type, 16#09#),
      11 => to_slv(opcode_type, 16#06#),
      12 => to_slv(opcode_type, 16#0F#),
      13 => to_slv(opcode_type, 16#0A#),
      14 => to_slv(opcode_type, 16#09#),
      15 => to_slv(opcode_type, 16#0B#),
      16 => to_slv(opcode_type, 16#0E#),
      17 => to_slv(opcode_type, 16#09#),
      18 => to_slv(opcode_type, 16#06#),
      19 => to_slv(opcode_type, 16#0D#),
      20 => to_slv(opcode_type, 16#0A#),
      21 => to_slv(opcode_type, 16#06#),
      22 => to_slv(opcode_type, 16#0B#),
      23 => to_slv(opcode_type, 16#10#),
      24 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#08#),
      33 => to_slv(opcode_type, 16#07#),
      34 => to_slv(opcode_type, 16#03#),
      35 => to_slv(opcode_type, 16#07#),
      36 => to_slv(opcode_type, 16#D8#),
      37 => to_slv(opcode_type, 16#0F#),
      38 => to_slv(opcode_type, 16#01#),
      39 => to_slv(opcode_type, 16#07#),
      40 => to_slv(opcode_type, 16#0B#),
      41 => to_slv(opcode_type, 16#0F#),
      42 => to_slv(opcode_type, 16#07#),
      43 => to_slv(opcode_type, 16#08#),
      44 => to_slv(opcode_type, 16#04#),
      45 => to_slv(opcode_type, 16#0A#),
      46 => to_slv(opcode_type, 16#06#),
      47 => to_slv(opcode_type, 16#0B#),
      48 => to_slv(opcode_type, 16#0A#),
      49 => to_slv(opcode_type, 16#08#),
      50 => to_slv(opcode_type, 16#07#),
      51 => to_slv(opcode_type, 16#0D#),
      52 => to_slv(opcode_type, 16#0B#),
      53 => to_slv(opcode_type, 16#06#),
      54 => to_slv(opcode_type, 16#0A#),
      55 => to_slv(opcode_type, 16#0C#),
      56 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#07#),
      65 => to_slv(opcode_type, 16#02#),
      66 => to_slv(opcode_type, 16#08#),
      67 => to_slv(opcode_type, 16#08#),
      68 => to_slv(opcode_type, 16#0A#),
      69 => to_slv(opcode_type, 16#0A#),
      70 => to_slv(opcode_type, 16#07#),
      71 => to_slv(opcode_type, 16#5B#),
      72 => to_slv(opcode_type, 16#0C#),
      73 => to_slv(opcode_type, 16#09#),
      74 => to_slv(opcode_type, 16#06#),
      75 => to_slv(opcode_type, 16#08#),
      76 => to_slv(opcode_type, 16#0D#),
      77 => to_slv(opcode_type, 16#0E#),
      78 => to_slv(opcode_type, 16#06#),
      79 => to_slv(opcode_type, 16#0E#),
      80 => to_slv(opcode_type, 16#11#),
      81 => to_slv(opcode_type, 16#08#),
      82 => to_slv(opcode_type, 16#06#),
      83 => to_slv(opcode_type, 16#0D#),
      84 => to_slv(opcode_type, 16#10#),
      85 => to_slv(opcode_type, 16#07#),
      86 => to_slv(opcode_type, 16#0F#),
      87 => to_slv(opcode_type, 16#0C#),
      88 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#08#),
      97 => to_slv(opcode_type, 16#04#),
      98 => to_slv(opcode_type, 16#09#),
      99 => to_slv(opcode_type, 16#08#),
      100 => to_slv(opcode_type, 16#0F#),
      101 => to_slv(opcode_type, 16#0C#),
      102 => to_slv(opcode_type, 16#07#),
      103 => to_slv(opcode_type, 16#0E#),
      104 => to_slv(opcode_type, 16#10#),
      105 => to_slv(opcode_type, 16#06#),
      106 => to_slv(opcode_type, 16#06#),
      107 => to_slv(opcode_type, 16#08#),
      108 => to_slv(opcode_type, 16#DA#),
      109 => to_slv(opcode_type, 16#0A#),
      110 => to_slv(opcode_type, 16#09#),
      111 => to_slv(opcode_type, 16#0F#),
      112 => to_slv(opcode_type, 16#0B#),
      113 => to_slv(opcode_type, 16#07#),
      114 => to_slv(opcode_type, 16#08#),
      115 => to_slv(opcode_type, 16#11#),
      116 => to_slv(opcode_type, 16#0A#),
      117 => to_slv(opcode_type, 16#08#),
      118 => to_slv(opcode_type, 16#0F#),
      119 => to_slv(opcode_type, 16#0C#),
      120 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#08#),
      129 => to_slv(opcode_type, 16#06#),
      130 => to_slv(opcode_type, 16#04#),
      131 => to_slv(opcode_type, 16#06#),
      132 => to_slv(opcode_type, 16#10#),
      133 => to_slv(opcode_type, 16#10#),
      134 => to_slv(opcode_type, 16#07#),
      135 => to_slv(opcode_type, 16#02#),
      136 => to_slv(opcode_type, 16#83#),
      137 => to_slv(opcode_type, 16#04#),
      138 => to_slv(opcode_type, 16#0F#),
      139 => to_slv(opcode_type, 16#08#),
      140 => to_slv(opcode_type, 16#09#),
      141 => to_slv(opcode_type, 16#04#),
      142 => to_slv(opcode_type, 16#48#),
      143 => to_slv(opcode_type, 16#01#),
      144 => to_slv(opcode_type, 16#0B#),
      145 => to_slv(opcode_type, 16#06#),
      146 => to_slv(opcode_type, 16#08#),
      147 => to_slv(opcode_type, 16#0F#),
      148 => to_slv(opcode_type, 16#0C#),
      149 => to_slv(opcode_type, 16#07#),
      150 => to_slv(opcode_type, 16#0F#),
      151 => to_slv(opcode_type, 16#0F#),
      152 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#06#),
      161 => to_slv(opcode_type, 16#04#),
      162 => to_slv(opcode_type, 16#08#),
      163 => to_slv(opcode_type, 16#06#),
      164 => to_slv(opcode_type, 16#0A#),
      165 => to_slv(opcode_type, 16#0C#),
      166 => to_slv(opcode_type, 16#08#),
      167 => to_slv(opcode_type, 16#0F#),
      168 => to_slv(opcode_type, 16#E0#),
      169 => to_slv(opcode_type, 16#06#),
      170 => to_slv(opcode_type, 16#06#),
      171 => to_slv(opcode_type, 16#08#),
      172 => to_slv(opcode_type, 16#0A#),
      173 => to_slv(opcode_type, 16#0F#),
      174 => to_slv(opcode_type, 16#06#),
      175 => to_slv(opcode_type, 16#0A#),
      176 => to_slv(opcode_type, 16#10#),
      177 => to_slv(opcode_type, 16#06#),
      178 => to_slv(opcode_type, 16#06#),
      179 => to_slv(opcode_type, 16#0F#),
      180 => to_slv(opcode_type, 16#11#),
      181 => to_slv(opcode_type, 16#09#),
      182 => to_slv(opcode_type, 16#0E#),
      183 => to_slv(opcode_type, 16#0E#),
      184 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#08#),
      193 => to_slv(opcode_type, 16#04#),
      194 => to_slv(opcode_type, 16#06#),
      195 => to_slv(opcode_type, 16#06#),
      196 => to_slv(opcode_type, 16#11#),
      197 => to_slv(opcode_type, 16#40#),
      198 => to_slv(opcode_type, 16#06#),
      199 => to_slv(opcode_type, 16#0C#),
      200 => to_slv(opcode_type, 16#0B#),
      201 => to_slv(opcode_type, 16#06#),
      202 => to_slv(opcode_type, 16#06#),
      203 => to_slv(opcode_type, 16#07#),
      204 => to_slv(opcode_type, 16#0E#),
      205 => to_slv(opcode_type, 16#0F#),
      206 => to_slv(opcode_type, 16#07#),
      207 => to_slv(opcode_type, 16#0D#),
      208 => to_slv(opcode_type, 16#11#),
      209 => to_slv(opcode_type, 16#08#),
      210 => to_slv(opcode_type, 16#07#),
      211 => to_slv(opcode_type, 16#0B#),
      212 => to_slv(opcode_type, 16#0A#),
      213 => to_slv(opcode_type, 16#06#),
      214 => to_slv(opcode_type, 16#5A#),
      215 => to_slv(opcode_type, 16#0B#),
      216 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#09#),
      225 => to_slv(opcode_type, 16#03#),
      226 => to_slv(opcode_type, 16#08#),
      227 => to_slv(opcode_type, 16#07#),
      228 => to_slv(opcode_type, 16#0C#),
      229 => to_slv(opcode_type, 16#0F#),
      230 => to_slv(opcode_type, 16#06#),
      231 => to_slv(opcode_type, 16#2D#),
      232 => to_slv(opcode_type, 16#0D#),
      233 => to_slv(opcode_type, 16#09#),
      234 => to_slv(opcode_type, 16#06#),
      235 => to_slv(opcode_type, 16#08#),
      236 => to_slv(opcode_type, 16#11#),
      237 => to_slv(opcode_type, 16#0E#),
      238 => to_slv(opcode_type, 16#09#),
      239 => to_slv(opcode_type, 16#0E#),
      240 => to_slv(opcode_type, 16#0F#),
      241 => to_slv(opcode_type, 16#06#),
      242 => to_slv(opcode_type, 16#08#),
      243 => to_slv(opcode_type, 16#0C#),
      244 => to_slv(opcode_type, 16#0C#),
      245 => to_slv(opcode_type, 16#06#),
      246 => to_slv(opcode_type, 16#0B#),
      247 => to_slv(opcode_type, 16#A5#),
      248 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#06#),
      257 => to_slv(opcode_type, 16#06#),
      258 => to_slv(opcode_type, 16#09#),
      259 => to_slv(opcode_type, 16#02#),
      260 => to_slv(opcode_type, 16#0F#),
      261 => to_slv(opcode_type, 16#01#),
      262 => to_slv(opcode_type, 16#32#),
      263 => to_slv(opcode_type, 16#03#),
      264 => to_slv(opcode_type, 16#08#),
      265 => to_slv(opcode_type, 16#0B#),
      266 => to_slv(opcode_type, 16#0E#),
      267 => to_slv(opcode_type, 16#07#),
      268 => to_slv(opcode_type, 16#07#),
      269 => to_slv(opcode_type, 16#06#),
      270 => to_slv(opcode_type, 16#B6#),
      271 => to_slv(opcode_type, 16#0C#),
      272 => to_slv(opcode_type, 16#05#),
      273 => to_slv(opcode_type, 16#0C#),
      274 => to_slv(opcode_type, 16#07#),
      275 => to_slv(opcode_type, 16#05#),
      276 => to_slv(opcode_type, 16#10#),
      277 => to_slv(opcode_type, 16#06#),
      278 => to_slv(opcode_type, 16#0E#),
      279 => to_slv(opcode_type, 16#10#),
      280 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#02#),
      290 => to_slv(opcode_type, 16#07#),
      291 => to_slv(opcode_type, 16#08#),
      292 => to_slv(opcode_type, 16#0A#),
      293 => to_slv(opcode_type, 16#0F#),
      294 => to_slv(opcode_type, 16#06#),
      295 => to_slv(opcode_type, 16#0D#),
      296 => to_slv(opcode_type, 16#0A#),
      297 => to_slv(opcode_type, 16#06#),
      298 => to_slv(opcode_type, 16#08#),
      299 => to_slv(opcode_type, 16#07#),
      300 => to_slv(opcode_type, 16#0F#),
      301 => to_slv(opcode_type, 16#7D#),
      302 => to_slv(opcode_type, 16#09#),
      303 => to_slv(opcode_type, 16#0A#),
      304 => to_slv(opcode_type, 16#11#),
      305 => to_slv(opcode_type, 16#08#),
      306 => to_slv(opcode_type, 16#09#),
      307 => to_slv(opcode_type, 16#0D#),
      308 => to_slv(opcode_type, 16#10#),
      309 => to_slv(opcode_type, 16#09#),
      310 => to_slv(opcode_type, 16#0B#),
      311 => to_slv(opcode_type, 16#72#),
      312 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#08#),
      321 => to_slv(opcode_type, 16#04#),
      322 => to_slv(opcode_type, 16#08#),
      323 => to_slv(opcode_type, 16#09#),
      324 => to_slv(opcode_type, 16#0C#),
      325 => to_slv(opcode_type, 16#0D#),
      326 => to_slv(opcode_type, 16#08#),
      327 => to_slv(opcode_type, 16#0D#),
      328 => to_slv(opcode_type, 16#0E#),
      329 => to_slv(opcode_type, 16#08#),
      330 => to_slv(opcode_type, 16#09#),
      331 => to_slv(opcode_type, 16#06#),
      332 => to_slv(opcode_type, 16#C0#),
      333 => to_slv(opcode_type, 16#0A#),
      334 => to_slv(opcode_type, 16#08#),
      335 => to_slv(opcode_type, 16#0E#),
      336 => to_slv(opcode_type, 16#0F#),
      337 => to_slv(opcode_type, 16#09#),
      338 => to_slv(opcode_type, 16#09#),
      339 => to_slv(opcode_type, 16#0A#),
      340 => to_slv(opcode_type, 16#0C#),
      341 => to_slv(opcode_type, 16#09#),
      342 => to_slv(opcode_type, 16#0E#),
      343 => to_slv(opcode_type, 16#0C#),
      344 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#09#),
      353 => to_slv(opcode_type, 16#06#),
      354 => to_slv(opcode_type, 16#05#),
      355 => to_slv(opcode_type, 16#07#),
      356 => to_slv(opcode_type, 16#0E#),
      357 => to_slv(opcode_type, 16#0C#),
      358 => to_slv(opcode_type, 16#07#),
      359 => to_slv(opcode_type, 16#05#),
      360 => to_slv(opcode_type, 16#0C#),
      361 => to_slv(opcode_type, 16#02#),
      362 => to_slv(opcode_type, 16#11#),
      363 => to_slv(opcode_type, 16#07#),
      364 => to_slv(opcode_type, 16#09#),
      365 => to_slv(opcode_type, 16#03#),
      366 => to_slv(opcode_type, 16#11#),
      367 => to_slv(opcode_type, 16#08#),
      368 => to_slv(opcode_type, 16#0C#),
      369 => to_slv(opcode_type, 16#0E#),
      370 => to_slv(opcode_type, 16#09#),
      371 => to_slv(opcode_type, 16#07#),
      372 => to_slv(opcode_type, 16#0B#),
      373 => to_slv(opcode_type, 16#10#),
      374 => to_slv(opcode_type, 16#03#),
      375 => to_slv(opcode_type, 16#0F#),
      376 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#08#),
      385 => to_slv(opcode_type, 16#02#),
      386 => to_slv(opcode_type, 16#07#),
      387 => to_slv(opcode_type, 16#08#),
      388 => to_slv(opcode_type, 16#10#),
      389 => to_slv(opcode_type, 16#10#),
      390 => to_slv(opcode_type, 16#08#),
      391 => to_slv(opcode_type, 16#11#),
      392 => to_slv(opcode_type, 16#0B#),
      393 => to_slv(opcode_type, 16#06#),
      394 => to_slv(opcode_type, 16#07#),
      395 => to_slv(opcode_type, 16#06#),
      396 => to_slv(opcode_type, 16#0A#),
      397 => to_slv(opcode_type, 16#0E#),
      398 => to_slv(opcode_type, 16#08#),
      399 => to_slv(opcode_type, 16#0C#),
      400 => to_slv(opcode_type, 16#0C#),
      401 => to_slv(opcode_type, 16#09#),
      402 => to_slv(opcode_type, 16#09#),
      403 => to_slv(opcode_type, 16#0B#),
      404 => to_slv(opcode_type, 16#0E#),
      405 => to_slv(opcode_type, 16#07#),
      406 => to_slv(opcode_type, 16#0B#),
      407 => to_slv(opcode_type, 16#0B#),
      408 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#07#),
      417 => to_slv(opcode_type, 16#09#),
      418 => to_slv(opcode_type, 16#09#),
      419 => to_slv(opcode_type, 16#06#),
      420 => to_slv(opcode_type, 16#0A#),
      421 => to_slv(opcode_type, 16#0E#),
      422 => to_slv(opcode_type, 16#02#),
      423 => to_slv(opcode_type, 16#0B#),
      424 => to_slv(opcode_type, 16#07#),
      425 => to_slv(opcode_type, 16#02#),
      426 => to_slv(opcode_type, 16#0C#),
      427 => to_slv(opcode_type, 16#09#),
      428 => to_slv(opcode_type, 16#0B#),
      429 => to_slv(opcode_type, 16#0F#),
      430 => to_slv(opcode_type, 16#07#),
      431 => to_slv(opcode_type, 16#08#),
      432 => to_slv(opcode_type, 16#08#),
      433 => to_slv(opcode_type, 16#0F#),
      434 => to_slv(opcode_type, 16#0B#),
      435 => to_slv(opcode_type, 16#03#),
      436 => to_slv(opcode_type, 16#0A#),
      437 => to_slv(opcode_type, 16#06#),
      438 => to_slv(opcode_type, 16#0F#),
      439 => to_slv(opcode_type, 16#10#),
      440 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#07#),
      449 => to_slv(opcode_type, 16#03#),
      450 => to_slv(opcode_type, 16#06#),
      451 => to_slv(opcode_type, 16#06#),
      452 => to_slv(opcode_type, 16#0B#),
      453 => to_slv(opcode_type, 16#0D#),
      454 => to_slv(opcode_type, 16#08#),
      455 => to_slv(opcode_type, 16#11#),
      456 => to_slv(opcode_type, 16#0B#),
      457 => to_slv(opcode_type, 16#06#),
      458 => to_slv(opcode_type, 16#06#),
      459 => to_slv(opcode_type, 16#06#),
      460 => to_slv(opcode_type, 16#5D#),
      461 => to_slv(opcode_type, 16#58#),
      462 => to_slv(opcode_type, 16#08#),
      463 => to_slv(opcode_type, 16#0E#),
      464 => to_slv(opcode_type, 16#10#),
      465 => to_slv(opcode_type, 16#09#),
      466 => to_slv(opcode_type, 16#06#),
      467 => to_slv(opcode_type, 16#0C#),
      468 => to_slv(opcode_type, 16#0E#),
      469 => to_slv(opcode_type, 16#07#),
      470 => to_slv(opcode_type, 16#0C#),
      471 => to_slv(opcode_type, 16#10#),
      472 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#06#),
      481 => to_slv(opcode_type, 16#09#),
      482 => to_slv(opcode_type, 16#08#),
      483 => to_slv(opcode_type, 16#08#),
      484 => to_slv(opcode_type, 16#0E#),
      485 => to_slv(opcode_type, 16#11#),
      486 => to_slv(opcode_type, 16#08#),
      487 => to_slv(opcode_type, 16#11#),
      488 => to_slv(opcode_type, 16#0E#),
      489 => to_slv(opcode_type, 16#03#),
      490 => to_slv(opcode_type, 16#05#),
      491 => to_slv(opcode_type, 16#0A#),
      492 => to_slv(opcode_type, 16#09#),
      493 => to_slv(opcode_type, 16#09#),
      494 => to_slv(opcode_type, 16#08#),
      495 => to_slv(opcode_type, 16#A8#),
      496 => to_slv(opcode_type, 16#0D#),
      497 => to_slv(opcode_type, 16#04#),
      498 => to_slv(opcode_type, 16#89#),
      499 => to_slv(opcode_type, 16#09#),
      500 => to_slv(opcode_type, 16#03#),
      501 => to_slv(opcode_type, 16#11#),
      502 => to_slv(opcode_type, 16#03#),
      503 => to_slv(opcode_type, 16#D9#),
      504 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#04#),
      514 => to_slv(opcode_type, 16#09#),
      515 => to_slv(opcode_type, 16#08#),
      516 => to_slv(opcode_type, 16#0A#),
      517 => to_slv(opcode_type, 16#0C#),
      518 => to_slv(opcode_type, 16#07#),
      519 => to_slv(opcode_type, 16#0E#),
      520 => to_slv(opcode_type, 16#10#),
      521 => to_slv(opcode_type, 16#08#),
      522 => to_slv(opcode_type, 16#08#),
      523 => to_slv(opcode_type, 16#09#),
      524 => to_slv(opcode_type, 16#0D#),
      525 => to_slv(opcode_type, 16#77#),
      526 => to_slv(opcode_type, 16#09#),
      527 => to_slv(opcode_type, 16#0D#),
      528 => to_slv(opcode_type, 16#0B#),
      529 => to_slv(opcode_type, 16#06#),
      530 => to_slv(opcode_type, 16#07#),
      531 => to_slv(opcode_type, 16#0B#),
      532 => to_slv(opcode_type, 16#1B#),
      533 => to_slv(opcode_type, 16#07#),
      534 => to_slv(opcode_type, 16#11#),
      535 => to_slv(opcode_type, 16#0D#),
      536 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#07#),
      545 => to_slv(opcode_type, 16#07#),
      546 => to_slv(opcode_type, 16#02#),
      547 => to_slv(opcode_type, 16#01#),
      548 => to_slv(opcode_type, 16#0C#),
      549 => to_slv(opcode_type, 16#01#),
      550 => to_slv(opcode_type, 16#06#),
      551 => to_slv(opcode_type, 16#CD#),
      552 => to_slv(opcode_type, 16#0C#),
      553 => to_slv(opcode_type, 16#09#),
      554 => to_slv(opcode_type, 16#07#),
      555 => to_slv(opcode_type, 16#07#),
      556 => to_slv(opcode_type, 16#0F#),
      557 => to_slv(opcode_type, 16#0C#),
      558 => to_slv(opcode_type, 16#09#),
      559 => to_slv(opcode_type, 16#0F#),
      560 => to_slv(opcode_type, 16#0C#),
      561 => to_slv(opcode_type, 16#08#),
      562 => to_slv(opcode_type, 16#07#),
      563 => to_slv(opcode_type, 16#11#),
      564 => to_slv(opcode_type, 16#0F#),
      565 => to_slv(opcode_type, 16#06#),
      566 => to_slv(opcode_type, 16#33#),
      567 => to_slv(opcode_type, 16#0C#),
      568 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#07#),
      577 => to_slv(opcode_type, 16#02#),
      578 => to_slv(opcode_type, 16#07#),
      579 => to_slv(opcode_type, 16#07#),
      580 => to_slv(opcode_type, 16#0B#),
      581 => to_slv(opcode_type, 16#0D#),
      582 => to_slv(opcode_type, 16#06#),
      583 => to_slv(opcode_type, 16#11#),
      584 => to_slv(opcode_type, 16#0C#),
      585 => to_slv(opcode_type, 16#06#),
      586 => to_slv(opcode_type, 16#09#),
      587 => to_slv(opcode_type, 16#08#),
      588 => to_slv(opcode_type, 16#11#),
      589 => to_slv(opcode_type, 16#2A#),
      590 => to_slv(opcode_type, 16#06#),
      591 => to_slv(opcode_type, 16#0F#),
      592 => to_slv(opcode_type, 16#0A#),
      593 => to_slv(opcode_type, 16#09#),
      594 => to_slv(opcode_type, 16#06#),
      595 => to_slv(opcode_type, 16#7A#),
      596 => to_slv(opcode_type, 16#0A#),
      597 => to_slv(opcode_type, 16#09#),
      598 => to_slv(opcode_type, 16#10#),
      599 => to_slv(opcode_type, 16#10#),
      600 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#07#),
      609 => to_slv(opcode_type, 16#08#),
      610 => to_slv(opcode_type, 16#09#),
      611 => to_slv(opcode_type, 16#04#),
      612 => to_slv(opcode_type, 16#0A#),
      613 => to_slv(opcode_type, 16#03#),
      614 => to_slv(opcode_type, 16#0C#),
      615 => to_slv(opcode_type, 16#05#),
      616 => to_slv(opcode_type, 16#08#),
      617 => to_slv(opcode_type, 16#0E#),
      618 => to_slv(opcode_type, 16#0B#),
      619 => to_slv(opcode_type, 16#08#),
      620 => to_slv(opcode_type, 16#08#),
      621 => to_slv(opcode_type, 16#04#),
      622 => to_slv(opcode_type, 16#0D#),
      623 => to_slv(opcode_type, 16#02#),
      624 => to_slv(opcode_type, 16#0D#),
      625 => to_slv(opcode_type, 16#09#),
      626 => to_slv(opcode_type, 16#07#),
      627 => to_slv(opcode_type, 16#0A#),
      628 => to_slv(opcode_type, 16#0C#),
      629 => to_slv(opcode_type, 16#07#),
      630 => to_slv(opcode_type, 16#0D#),
      631 => to_slv(opcode_type, 16#0E#),
      632 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#09#),
      641 => to_slv(opcode_type, 16#02#),
      642 => to_slv(opcode_type, 16#07#),
      643 => to_slv(opcode_type, 16#06#),
      644 => to_slv(opcode_type, 16#0B#),
      645 => to_slv(opcode_type, 16#0F#),
      646 => to_slv(opcode_type, 16#07#),
      647 => to_slv(opcode_type, 16#11#),
      648 => to_slv(opcode_type, 16#0B#),
      649 => to_slv(opcode_type, 16#06#),
      650 => to_slv(opcode_type, 16#07#),
      651 => to_slv(opcode_type, 16#07#),
      652 => to_slv(opcode_type, 16#0C#),
      653 => to_slv(opcode_type, 16#A0#),
      654 => to_slv(opcode_type, 16#08#),
      655 => to_slv(opcode_type, 16#0A#),
      656 => to_slv(opcode_type, 16#A6#),
      657 => to_slv(opcode_type, 16#09#),
      658 => to_slv(opcode_type, 16#07#),
      659 => to_slv(opcode_type, 16#0A#),
      660 => to_slv(opcode_type, 16#0F#),
      661 => to_slv(opcode_type, 16#07#),
      662 => to_slv(opcode_type, 16#0C#),
      663 => to_slv(opcode_type, 16#0F#),
      664 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#09#),
      673 => to_slv(opcode_type, 16#09#),
      674 => to_slv(opcode_type, 16#03#),
      675 => to_slv(opcode_type, 16#06#),
      676 => to_slv(opcode_type, 16#11#),
      677 => to_slv(opcode_type, 16#0F#),
      678 => to_slv(opcode_type, 16#01#),
      679 => to_slv(opcode_type, 16#07#),
      680 => to_slv(opcode_type, 16#0D#),
      681 => to_slv(opcode_type, 16#0E#),
      682 => to_slv(opcode_type, 16#07#),
      683 => to_slv(opcode_type, 16#08#),
      684 => to_slv(opcode_type, 16#08#),
      685 => to_slv(opcode_type, 16#0F#),
      686 => to_slv(opcode_type, 16#0B#),
      687 => to_slv(opcode_type, 16#03#),
      688 => to_slv(opcode_type, 16#11#),
      689 => to_slv(opcode_type, 16#06#),
      690 => to_slv(opcode_type, 16#06#),
      691 => to_slv(opcode_type, 16#10#),
      692 => to_slv(opcode_type, 16#0F#),
      693 => to_slv(opcode_type, 16#09#),
      694 => to_slv(opcode_type, 16#0C#),
      695 => to_slv(opcode_type, 16#0F#),
      696 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#09#),
      705 => to_slv(opcode_type, 16#04#),
      706 => to_slv(opcode_type, 16#09#),
      707 => to_slv(opcode_type, 16#07#),
      708 => to_slv(opcode_type, 16#11#),
      709 => to_slv(opcode_type, 16#0A#),
      710 => to_slv(opcode_type, 16#08#),
      711 => to_slv(opcode_type, 16#0C#),
      712 => to_slv(opcode_type, 16#0A#),
      713 => to_slv(opcode_type, 16#08#),
      714 => to_slv(opcode_type, 16#08#),
      715 => to_slv(opcode_type, 16#08#),
      716 => to_slv(opcode_type, 16#0F#),
      717 => to_slv(opcode_type, 16#0B#),
      718 => to_slv(opcode_type, 16#07#),
      719 => to_slv(opcode_type, 16#0E#),
      720 => to_slv(opcode_type, 16#0A#),
      721 => to_slv(opcode_type, 16#09#),
      722 => to_slv(opcode_type, 16#06#),
      723 => to_slv(opcode_type, 16#0F#),
      724 => to_slv(opcode_type, 16#0C#),
      725 => to_slv(opcode_type, 16#08#),
      726 => to_slv(opcode_type, 16#0A#),
      727 => to_slv(opcode_type, 16#10#),
      728 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#07#),
      737 => to_slv(opcode_type, 16#01#),
      738 => to_slv(opcode_type, 16#06#),
      739 => to_slv(opcode_type, 16#09#),
      740 => to_slv(opcode_type, 16#0A#),
      741 => to_slv(opcode_type, 16#0C#),
      742 => to_slv(opcode_type, 16#08#),
      743 => to_slv(opcode_type, 16#75#),
      744 => to_slv(opcode_type, 16#0D#),
      745 => to_slv(opcode_type, 16#09#),
      746 => to_slv(opcode_type, 16#07#),
      747 => to_slv(opcode_type, 16#09#),
      748 => to_slv(opcode_type, 16#11#),
      749 => to_slv(opcode_type, 16#0C#),
      750 => to_slv(opcode_type, 16#06#),
      751 => to_slv(opcode_type, 16#0E#),
      752 => to_slv(opcode_type, 16#0D#),
      753 => to_slv(opcode_type, 16#06#),
      754 => to_slv(opcode_type, 16#09#),
      755 => to_slv(opcode_type, 16#0F#),
      756 => to_slv(opcode_type, 16#0B#),
      757 => to_slv(opcode_type, 16#09#),
      758 => to_slv(opcode_type, 16#0B#),
      759 => to_slv(opcode_type, 16#0F#),
      760 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#07#),
      769 => to_slv(opcode_type, 16#03#),
      770 => to_slv(opcode_type, 16#06#),
      771 => to_slv(opcode_type, 16#08#),
      772 => to_slv(opcode_type, 16#0A#),
      773 => to_slv(opcode_type, 16#10#),
      774 => to_slv(opcode_type, 16#09#),
      775 => to_slv(opcode_type, 16#10#),
      776 => to_slv(opcode_type, 16#0A#),
      777 => to_slv(opcode_type, 16#06#),
      778 => to_slv(opcode_type, 16#09#),
      779 => to_slv(opcode_type, 16#06#),
      780 => to_slv(opcode_type, 16#10#),
      781 => to_slv(opcode_type, 16#0B#),
      782 => to_slv(opcode_type, 16#06#),
      783 => to_slv(opcode_type, 16#0A#),
      784 => to_slv(opcode_type, 16#0A#),
      785 => to_slv(opcode_type, 16#08#),
      786 => to_slv(opcode_type, 16#06#),
      787 => to_slv(opcode_type, 16#11#),
      788 => to_slv(opcode_type, 16#0F#),
      789 => to_slv(opcode_type, 16#07#),
      790 => to_slv(opcode_type, 16#0B#),
      791 => to_slv(opcode_type, 16#0C#),
      792 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#07#),
      801 => to_slv(opcode_type, 16#06#),
      802 => to_slv(opcode_type, 16#07#),
      803 => to_slv(opcode_type, 16#01#),
      804 => to_slv(opcode_type, 16#11#),
      805 => to_slv(opcode_type, 16#07#),
      806 => to_slv(opcode_type, 16#0C#),
      807 => to_slv(opcode_type, 16#0B#),
      808 => to_slv(opcode_type, 16#08#),
      809 => to_slv(opcode_type, 16#04#),
      810 => to_slv(opcode_type, 16#0C#),
      811 => to_slv(opcode_type, 16#01#),
      812 => to_slv(opcode_type, 16#11#),
      813 => to_slv(opcode_type, 16#08#),
      814 => to_slv(opcode_type, 16#05#),
      815 => to_slv(opcode_type, 16#07#),
      816 => to_slv(opcode_type, 16#11#),
      817 => to_slv(opcode_type, 16#11#),
      818 => to_slv(opcode_type, 16#09#),
      819 => to_slv(opcode_type, 16#01#),
      820 => to_slv(opcode_type, 16#0C#),
      821 => to_slv(opcode_type, 16#07#),
      822 => to_slv(opcode_type, 16#0E#),
      823 => to_slv(opcode_type, 16#0C#),
      824 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#06#),
      833 => to_slv(opcode_type, 16#06#),
      834 => to_slv(opcode_type, 16#07#),
      835 => to_slv(opcode_type, 16#04#),
      836 => to_slv(opcode_type, 16#0F#),
      837 => to_slv(opcode_type, 16#04#),
      838 => to_slv(opcode_type, 16#10#),
      839 => to_slv(opcode_type, 16#05#),
      840 => to_slv(opcode_type, 16#04#),
      841 => to_slv(opcode_type, 16#0E#),
      842 => to_slv(opcode_type, 16#09#),
      843 => to_slv(opcode_type, 16#06#),
      844 => to_slv(opcode_type, 16#04#),
      845 => to_slv(opcode_type, 16#28#),
      846 => to_slv(opcode_type, 16#06#),
      847 => to_slv(opcode_type, 16#0F#),
      848 => to_slv(opcode_type, 16#10#),
      849 => to_slv(opcode_type, 16#07#),
      850 => to_slv(opcode_type, 16#06#),
      851 => to_slv(opcode_type, 16#0C#),
      852 => to_slv(opcode_type, 16#0A#),
      853 => to_slv(opcode_type, 16#06#),
      854 => to_slv(opcode_type, 16#0A#),
      855 => to_slv(opcode_type, 16#0B#),
      856 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#08#),
      865 => to_slv(opcode_type, 16#03#),
      866 => to_slv(opcode_type, 16#06#),
      867 => to_slv(opcode_type, 16#09#),
      868 => to_slv(opcode_type, 16#0E#),
      869 => to_slv(opcode_type, 16#60#),
      870 => to_slv(opcode_type, 16#07#),
      871 => to_slv(opcode_type, 16#10#),
      872 => to_slv(opcode_type, 16#10#),
      873 => to_slv(opcode_type, 16#07#),
      874 => to_slv(opcode_type, 16#07#),
      875 => to_slv(opcode_type, 16#09#),
      876 => to_slv(opcode_type, 16#10#),
      877 => to_slv(opcode_type, 16#0A#),
      878 => to_slv(opcode_type, 16#09#),
      879 => to_slv(opcode_type, 16#11#),
      880 => to_slv(opcode_type, 16#0F#),
      881 => to_slv(opcode_type, 16#07#),
      882 => to_slv(opcode_type, 16#09#),
      883 => to_slv(opcode_type, 16#0E#),
      884 => to_slv(opcode_type, 16#12#),
      885 => to_slv(opcode_type, 16#06#),
      886 => to_slv(opcode_type, 16#0A#),
      887 => to_slv(opcode_type, 16#0F#),
      888 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#08#),
      897 => to_slv(opcode_type, 16#06#),
      898 => to_slv(opcode_type, 16#08#),
      899 => to_slv(opcode_type, 16#05#),
      900 => to_slv(opcode_type, 16#0B#),
      901 => to_slv(opcode_type, 16#07#),
      902 => to_slv(opcode_type, 16#0B#),
      903 => to_slv(opcode_type, 16#11#),
      904 => to_slv(opcode_type, 16#05#),
      905 => to_slv(opcode_type, 16#01#),
      906 => to_slv(opcode_type, 16#0B#),
      907 => to_slv(opcode_type, 16#06#),
      908 => to_slv(opcode_type, 16#09#),
      909 => to_slv(opcode_type, 16#04#),
      910 => to_slv(opcode_type, 16#A6#),
      911 => to_slv(opcode_type, 16#01#),
      912 => to_slv(opcode_type, 16#5D#),
      913 => to_slv(opcode_type, 16#09#),
      914 => to_slv(opcode_type, 16#06#),
      915 => to_slv(opcode_type, 16#0B#),
      916 => to_slv(opcode_type, 16#0A#),
      917 => to_slv(opcode_type, 16#06#),
      918 => to_slv(opcode_type, 16#0A#),
      919 => to_slv(opcode_type, 16#11#),
      920 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#07#),
      929 => to_slv(opcode_type, 16#05#),
      930 => to_slv(opcode_type, 16#06#),
      931 => to_slv(opcode_type, 16#06#),
      932 => to_slv(opcode_type, 16#12#),
      933 => to_slv(opcode_type, 16#0A#),
      934 => to_slv(opcode_type, 16#07#),
      935 => to_slv(opcode_type, 16#0A#),
      936 => to_slv(opcode_type, 16#0C#),
      937 => to_slv(opcode_type, 16#09#),
      938 => to_slv(opcode_type, 16#08#),
      939 => to_slv(opcode_type, 16#07#),
      940 => to_slv(opcode_type, 16#10#),
      941 => to_slv(opcode_type, 16#0A#),
      942 => to_slv(opcode_type, 16#06#),
      943 => to_slv(opcode_type, 16#10#),
      944 => to_slv(opcode_type, 16#0B#),
      945 => to_slv(opcode_type, 16#08#),
      946 => to_slv(opcode_type, 16#08#),
      947 => to_slv(opcode_type, 16#0D#),
      948 => to_slv(opcode_type, 16#0A#),
      949 => to_slv(opcode_type, 16#09#),
      950 => to_slv(opcode_type, 16#0C#),
      951 => to_slv(opcode_type, 16#0F#),
      952 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#06#),
      961 => to_slv(opcode_type, 16#05#),
      962 => to_slv(opcode_type, 16#08#),
      963 => to_slv(opcode_type, 16#07#),
      964 => to_slv(opcode_type, 16#59#),
      965 => to_slv(opcode_type, 16#0C#),
      966 => to_slv(opcode_type, 16#09#),
      967 => to_slv(opcode_type, 16#0C#),
      968 => to_slv(opcode_type, 16#10#),
      969 => to_slv(opcode_type, 16#08#),
      970 => to_slv(opcode_type, 16#08#),
      971 => to_slv(opcode_type, 16#08#),
      972 => to_slv(opcode_type, 16#0A#),
      973 => to_slv(opcode_type, 16#0B#),
      974 => to_slv(opcode_type, 16#06#),
      975 => to_slv(opcode_type, 16#0F#),
      976 => to_slv(opcode_type, 16#0B#),
      977 => to_slv(opcode_type, 16#07#),
      978 => to_slv(opcode_type, 16#07#),
      979 => to_slv(opcode_type, 16#11#),
      980 => to_slv(opcode_type, 16#9B#),
      981 => to_slv(opcode_type, 16#07#),
      982 => to_slv(opcode_type, 16#0F#),
      983 => to_slv(opcode_type, 16#11#),
      984 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#07#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#08#),
      995 => to_slv(opcode_type, 16#03#),
      996 => to_slv(opcode_type, 16#10#),
      997 => to_slv(opcode_type, 16#06#),
      998 => to_slv(opcode_type, 16#0D#),
      999 => to_slv(opcode_type, 16#63#),
      1000 => to_slv(opcode_type, 16#01#),
      1001 => to_slv(opcode_type, 16#03#),
      1002 => to_slv(opcode_type, 16#0D#),
      1003 => to_slv(opcode_type, 16#06#),
      1004 => to_slv(opcode_type, 16#08#),
      1005 => to_slv(opcode_type, 16#08#),
      1006 => to_slv(opcode_type, 16#0A#),
      1007 => to_slv(opcode_type, 16#10#),
      1008 => to_slv(opcode_type, 16#01#),
      1009 => to_slv(opcode_type, 16#10#),
      1010 => to_slv(opcode_type, 16#08#),
      1011 => to_slv(opcode_type, 16#01#),
      1012 => to_slv(opcode_type, 16#0D#),
      1013 => to_slv(opcode_type, 16#09#),
      1014 => to_slv(opcode_type, 16#0E#),
      1015 => to_slv(opcode_type, 16#0A#),
      1016 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#08#),
      1025 => to_slv(opcode_type, 16#05#),
      1026 => to_slv(opcode_type, 16#09#),
      1027 => to_slv(opcode_type, 16#06#),
      1028 => to_slv(opcode_type, 16#0D#),
      1029 => to_slv(opcode_type, 16#0D#),
      1030 => to_slv(opcode_type, 16#06#),
      1031 => to_slv(opcode_type, 16#0E#),
      1032 => to_slv(opcode_type, 16#11#),
      1033 => to_slv(opcode_type, 16#06#),
      1034 => to_slv(opcode_type, 16#06#),
      1035 => to_slv(opcode_type, 16#09#),
      1036 => to_slv(opcode_type, 16#0D#),
      1037 => to_slv(opcode_type, 16#0A#),
      1038 => to_slv(opcode_type, 16#06#),
      1039 => to_slv(opcode_type, 16#0E#),
      1040 => to_slv(opcode_type, 16#11#),
      1041 => to_slv(opcode_type, 16#07#),
      1042 => to_slv(opcode_type, 16#08#),
      1043 => to_slv(opcode_type, 16#83#),
      1044 => to_slv(opcode_type, 16#0D#),
      1045 => to_slv(opcode_type, 16#08#),
      1046 => to_slv(opcode_type, 16#0C#),
      1047 => to_slv(opcode_type, 16#10#),
      1048 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#09#),
      1057 => to_slv(opcode_type, 16#02#),
      1058 => to_slv(opcode_type, 16#07#),
      1059 => to_slv(opcode_type, 16#09#),
      1060 => to_slv(opcode_type, 16#0B#),
      1061 => to_slv(opcode_type, 16#0D#),
      1062 => to_slv(opcode_type, 16#09#),
      1063 => to_slv(opcode_type, 16#0E#),
      1064 => to_slv(opcode_type, 16#10#),
      1065 => to_slv(opcode_type, 16#08#),
      1066 => to_slv(opcode_type, 16#08#),
      1067 => to_slv(opcode_type, 16#06#),
      1068 => to_slv(opcode_type, 16#11#),
      1069 => to_slv(opcode_type, 16#11#),
      1070 => to_slv(opcode_type, 16#08#),
      1071 => to_slv(opcode_type, 16#0E#),
      1072 => to_slv(opcode_type, 16#0F#),
      1073 => to_slv(opcode_type, 16#08#),
      1074 => to_slv(opcode_type, 16#09#),
      1075 => to_slv(opcode_type, 16#0E#),
      1076 => to_slv(opcode_type, 16#0A#),
      1077 => to_slv(opcode_type, 16#09#),
      1078 => to_slv(opcode_type, 16#0E#),
      1079 => to_slv(opcode_type, 16#10#),
      1080 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#08#),
      1089 => to_slv(opcode_type, 16#03#),
      1090 => to_slv(opcode_type, 16#09#),
      1091 => to_slv(opcode_type, 16#09#),
      1092 => to_slv(opcode_type, 16#0D#),
      1093 => to_slv(opcode_type, 16#0C#),
      1094 => to_slv(opcode_type, 16#07#),
      1095 => to_slv(opcode_type, 16#11#),
      1096 => to_slv(opcode_type, 16#E3#),
      1097 => to_slv(opcode_type, 16#09#),
      1098 => to_slv(opcode_type, 16#08#),
      1099 => to_slv(opcode_type, 16#08#),
      1100 => to_slv(opcode_type, 16#0E#),
      1101 => to_slv(opcode_type, 16#11#),
      1102 => to_slv(opcode_type, 16#06#),
      1103 => to_slv(opcode_type, 16#30#),
      1104 => to_slv(opcode_type, 16#11#),
      1105 => to_slv(opcode_type, 16#08#),
      1106 => to_slv(opcode_type, 16#07#),
      1107 => to_slv(opcode_type, 16#10#),
      1108 => to_slv(opcode_type, 16#0A#),
      1109 => to_slv(opcode_type, 16#06#),
      1110 => to_slv(opcode_type, 16#0F#),
      1111 => to_slv(opcode_type, 16#0F#),
      1112 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#09#),
      1121 => to_slv(opcode_type, 16#06#),
      1122 => to_slv(opcode_type, 16#02#),
      1123 => to_slv(opcode_type, 16#07#),
      1124 => to_slv(opcode_type, 16#0E#),
      1125 => to_slv(opcode_type, 16#0B#),
      1126 => to_slv(opcode_type, 16#08#),
      1127 => to_slv(opcode_type, 16#06#),
      1128 => to_slv(opcode_type, 16#0C#),
      1129 => to_slv(opcode_type, 16#0F#),
      1130 => to_slv(opcode_type, 16#08#),
      1131 => to_slv(opcode_type, 16#11#),
      1132 => to_slv(opcode_type, 16#0B#),
      1133 => to_slv(opcode_type, 16#07#),
      1134 => to_slv(opcode_type, 16#01#),
      1135 => to_slv(opcode_type, 16#02#),
      1136 => to_slv(opcode_type, 16#0A#),
      1137 => to_slv(opcode_type, 16#06#),
      1138 => to_slv(opcode_type, 16#08#),
      1139 => to_slv(opcode_type, 16#11#),
      1140 => to_slv(opcode_type, 16#0F#),
      1141 => to_slv(opcode_type, 16#07#),
      1142 => to_slv(opcode_type, 16#0B#),
      1143 => to_slv(opcode_type, 16#0B#),
      1144 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#07#),
      1153 => to_slv(opcode_type, 16#08#),
      1154 => to_slv(opcode_type, 16#03#),
      1155 => to_slv(opcode_type, 16#06#),
      1156 => to_slv(opcode_type, 16#11#),
      1157 => to_slv(opcode_type, 16#32#),
      1158 => to_slv(opcode_type, 16#04#),
      1159 => to_slv(opcode_type, 16#08#),
      1160 => to_slv(opcode_type, 16#0E#),
      1161 => to_slv(opcode_type, 16#10#),
      1162 => to_slv(opcode_type, 16#08#),
      1163 => to_slv(opcode_type, 16#06#),
      1164 => to_slv(opcode_type, 16#01#),
      1165 => to_slv(opcode_type, 16#0E#),
      1166 => to_slv(opcode_type, 16#08#),
      1167 => to_slv(opcode_type, 16#7E#),
      1168 => to_slv(opcode_type, 16#0E#),
      1169 => to_slv(opcode_type, 16#07#),
      1170 => to_slv(opcode_type, 16#07#),
      1171 => to_slv(opcode_type, 16#10#),
      1172 => to_slv(opcode_type, 16#0D#),
      1173 => to_slv(opcode_type, 16#08#),
      1174 => to_slv(opcode_type, 16#0F#),
      1175 => to_slv(opcode_type, 16#10#),
      1176 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#08#),
      1185 => to_slv(opcode_type, 16#01#),
      1186 => to_slv(opcode_type, 16#06#),
      1187 => to_slv(opcode_type, 16#08#),
      1188 => to_slv(opcode_type, 16#0B#),
      1189 => to_slv(opcode_type, 16#10#),
      1190 => to_slv(opcode_type, 16#07#),
      1191 => to_slv(opcode_type, 16#0C#),
      1192 => to_slv(opcode_type, 16#10#),
      1193 => to_slv(opcode_type, 16#09#),
      1194 => to_slv(opcode_type, 16#09#),
      1195 => to_slv(opcode_type, 16#09#),
      1196 => to_slv(opcode_type, 16#0C#),
      1197 => to_slv(opcode_type, 16#0A#),
      1198 => to_slv(opcode_type, 16#07#),
      1199 => to_slv(opcode_type, 16#0A#),
      1200 => to_slv(opcode_type, 16#10#),
      1201 => to_slv(opcode_type, 16#08#),
      1202 => to_slv(opcode_type, 16#07#),
      1203 => to_slv(opcode_type, 16#D8#),
      1204 => to_slv(opcode_type, 16#0B#),
      1205 => to_slv(opcode_type, 16#08#),
      1206 => to_slv(opcode_type, 16#0C#),
      1207 => to_slv(opcode_type, 16#0E#),
      1208 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#06#),
      1217 => to_slv(opcode_type, 16#08#),
      1218 => to_slv(opcode_type, 16#02#),
      1219 => to_slv(opcode_type, 16#05#),
      1220 => to_slv(opcode_type, 16#0A#),
      1221 => to_slv(opcode_type, 16#01#),
      1222 => to_slv(opcode_type, 16#09#),
      1223 => to_slv(opcode_type, 16#0F#),
      1224 => to_slv(opcode_type, 16#0A#),
      1225 => to_slv(opcode_type, 16#09#),
      1226 => to_slv(opcode_type, 16#06#),
      1227 => to_slv(opcode_type, 16#06#),
      1228 => to_slv(opcode_type, 16#10#),
      1229 => to_slv(opcode_type, 16#0E#),
      1230 => to_slv(opcode_type, 16#07#),
      1231 => to_slv(opcode_type, 16#DC#),
      1232 => to_slv(opcode_type, 16#0B#),
      1233 => to_slv(opcode_type, 16#06#),
      1234 => to_slv(opcode_type, 16#07#),
      1235 => to_slv(opcode_type, 16#0D#),
      1236 => to_slv(opcode_type, 16#0B#),
      1237 => to_slv(opcode_type, 16#06#),
      1238 => to_slv(opcode_type, 16#10#),
      1239 => to_slv(opcode_type, 16#C6#),
      1240 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#07#),
      1249 => to_slv(opcode_type, 16#07#),
      1250 => to_slv(opcode_type, 16#06#),
      1251 => to_slv(opcode_type, 16#01#),
      1252 => to_slv(opcode_type, 16#0D#),
      1253 => to_slv(opcode_type, 16#03#),
      1254 => to_slv(opcode_type, 16#11#),
      1255 => to_slv(opcode_type, 16#04#),
      1256 => to_slv(opcode_type, 16#02#),
      1257 => to_slv(opcode_type, 16#11#),
      1258 => to_slv(opcode_type, 16#08#),
      1259 => to_slv(opcode_type, 16#07#),
      1260 => to_slv(opcode_type, 16#06#),
      1261 => to_slv(opcode_type, 16#0D#),
      1262 => to_slv(opcode_type, 16#0A#),
      1263 => to_slv(opcode_type, 16#01#),
      1264 => to_slv(opcode_type, 16#11#),
      1265 => to_slv(opcode_type, 16#06#),
      1266 => to_slv(opcode_type, 16#09#),
      1267 => to_slv(opcode_type, 16#11#),
      1268 => to_slv(opcode_type, 16#11#),
      1269 => to_slv(opcode_type, 16#06#),
      1270 => to_slv(opcode_type, 16#0F#),
      1271 => to_slv(opcode_type, 16#0F#),
      1272 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#08#),
      1282 => to_slv(opcode_type, 16#01#),
      1283 => to_slv(opcode_type, 16#02#),
      1284 => to_slv(opcode_type, 16#8E#),
      1285 => to_slv(opcode_type, 16#05#),
      1286 => to_slv(opcode_type, 16#08#),
      1287 => to_slv(opcode_type, 16#11#),
      1288 => to_slv(opcode_type, 16#0D#),
      1289 => to_slv(opcode_type, 16#09#),
      1290 => to_slv(opcode_type, 16#09#),
      1291 => to_slv(opcode_type, 16#07#),
      1292 => to_slv(opcode_type, 16#10#),
      1293 => to_slv(opcode_type, 16#11#),
      1294 => to_slv(opcode_type, 16#06#),
      1295 => to_slv(opcode_type, 16#0F#),
      1296 => to_slv(opcode_type, 16#0B#),
      1297 => to_slv(opcode_type, 16#07#),
      1298 => to_slv(opcode_type, 16#07#),
      1299 => to_slv(opcode_type, 16#3A#),
      1300 => to_slv(opcode_type, 16#0F#),
      1301 => to_slv(opcode_type, 16#09#),
      1302 => to_slv(opcode_type, 16#0B#),
      1303 => to_slv(opcode_type, 16#27#),
      1304 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#08#),
      1313 => to_slv(opcode_type, 16#07#),
      1314 => to_slv(opcode_type, 16#04#),
      1315 => to_slv(opcode_type, 16#01#),
      1316 => to_slv(opcode_type, 16#11#),
      1317 => to_slv(opcode_type, 16#03#),
      1318 => to_slv(opcode_type, 16#08#),
      1319 => to_slv(opcode_type, 16#0D#),
      1320 => to_slv(opcode_type, 16#0F#),
      1321 => to_slv(opcode_type, 16#09#),
      1322 => to_slv(opcode_type, 16#08#),
      1323 => to_slv(opcode_type, 16#09#),
      1324 => to_slv(opcode_type, 16#0E#),
      1325 => to_slv(opcode_type, 16#0D#),
      1326 => to_slv(opcode_type, 16#08#),
      1327 => to_slv(opcode_type, 16#0D#),
      1328 => to_slv(opcode_type, 16#0B#),
      1329 => to_slv(opcode_type, 16#09#),
      1330 => to_slv(opcode_type, 16#07#),
      1331 => to_slv(opcode_type, 16#0E#),
      1332 => to_slv(opcode_type, 16#0D#),
      1333 => to_slv(opcode_type, 16#06#),
      1334 => to_slv(opcode_type, 16#10#),
      1335 => to_slv(opcode_type, 16#0A#),
      1336 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#08#),
      1345 => to_slv(opcode_type, 16#08#),
      1346 => to_slv(opcode_type, 16#04#),
      1347 => to_slv(opcode_type, 16#04#),
      1348 => to_slv(opcode_type, 16#0D#),
      1349 => to_slv(opcode_type, 16#01#),
      1350 => to_slv(opcode_type, 16#06#),
      1351 => to_slv(opcode_type, 16#0C#),
      1352 => to_slv(opcode_type, 16#0E#),
      1353 => to_slv(opcode_type, 16#06#),
      1354 => to_slv(opcode_type, 16#07#),
      1355 => to_slv(opcode_type, 16#09#),
      1356 => to_slv(opcode_type, 16#0B#),
      1357 => to_slv(opcode_type, 16#0E#),
      1358 => to_slv(opcode_type, 16#07#),
      1359 => to_slv(opcode_type, 16#0B#),
      1360 => to_slv(opcode_type, 16#0E#),
      1361 => to_slv(opcode_type, 16#07#),
      1362 => to_slv(opcode_type, 16#06#),
      1363 => to_slv(opcode_type, 16#10#),
      1364 => to_slv(opcode_type, 16#10#),
      1365 => to_slv(opcode_type, 16#08#),
      1366 => to_slv(opcode_type, 16#0D#),
      1367 => to_slv(opcode_type, 16#66#),
      1368 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#07#),
      1377 => to_slv(opcode_type, 16#01#),
      1378 => to_slv(opcode_type, 16#07#),
      1379 => to_slv(opcode_type, 16#08#),
      1380 => to_slv(opcode_type, 16#0C#),
      1381 => to_slv(opcode_type, 16#0F#),
      1382 => to_slv(opcode_type, 16#06#),
      1383 => to_slv(opcode_type, 16#0B#),
      1384 => to_slv(opcode_type, 16#0D#),
      1385 => to_slv(opcode_type, 16#06#),
      1386 => to_slv(opcode_type, 16#08#),
      1387 => to_slv(opcode_type, 16#06#),
      1388 => to_slv(opcode_type, 16#0F#),
      1389 => to_slv(opcode_type, 16#0E#),
      1390 => to_slv(opcode_type, 16#08#),
      1391 => to_slv(opcode_type, 16#10#),
      1392 => to_slv(opcode_type, 16#0A#),
      1393 => to_slv(opcode_type, 16#07#),
      1394 => to_slv(opcode_type, 16#08#),
      1395 => to_slv(opcode_type, 16#8E#),
      1396 => to_slv(opcode_type, 16#8B#),
      1397 => to_slv(opcode_type, 16#09#),
      1398 => to_slv(opcode_type, 16#DC#),
      1399 => to_slv(opcode_type, 16#0B#),
      1400 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#08#),
      1409 => to_slv(opcode_type, 16#09#),
      1410 => to_slv(opcode_type, 16#02#),
      1411 => to_slv(opcode_type, 16#06#),
      1412 => to_slv(opcode_type, 16#0E#),
      1413 => to_slv(opcode_type, 16#10#),
      1414 => to_slv(opcode_type, 16#08#),
      1415 => to_slv(opcode_type, 16#02#),
      1416 => to_slv(opcode_type, 16#0B#),
      1417 => to_slv(opcode_type, 16#08#),
      1418 => to_slv(opcode_type, 16#11#),
      1419 => to_slv(opcode_type, 16#0D#),
      1420 => to_slv(opcode_type, 16#07#),
      1421 => to_slv(opcode_type, 16#06#),
      1422 => to_slv(opcode_type, 16#03#),
      1423 => to_slv(opcode_type, 16#0C#),
      1424 => to_slv(opcode_type, 16#06#),
      1425 => to_slv(opcode_type, 16#0F#),
      1426 => to_slv(opcode_type, 16#11#),
      1427 => to_slv(opcode_type, 16#07#),
      1428 => to_slv(opcode_type, 16#07#),
      1429 => to_slv(opcode_type, 16#0B#),
      1430 => to_slv(opcode_type, 16#0B#),
      1431 => to_slv(opcode_type, 16#10#),
      1432 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#06#),
      1441 => to_slv(opcode_type, 16#05#),
      1442 => to_slv(opcode_type, 16#09#),
      1443 => to_slv(opcode_type, 16#08#),
      1444 => to_slv(opcode_type, 16#BD#),
      1445 => to_slv(opcode_type, 16#0A#),
      1446 => to_slv(opcode_type, 16#08#),
      1447 => to_slv(opcode_type, 16#0F#),
      1448 => to_slv(opcode_type, 16#0A#),
      1449 => to_slv(opcode_type, 16#08#),
      1450 => to_slv(opcode_type, 16#09#),
      1451 => to_slv(opcode_type, 16#08#),
      1452 => to_slv(opcode_type, 16#0D#),
      1453 => to_slv(opcode_type, 16#0C#),
      1454 => to_slv(opcode_type, 16#07#),
      1455 => to_slv(opcode_type, 16#0F#),
      1456 => to_slv(opcode_type, 16#11#),
      1457 => to_slv(opcode_type, 16#09#),
      1458 => to_slv(opcode_type, 16#06#),
      1459 => to_slv(opcode_type, 16#0F#),
      1460 => to_slv(opcode_type, 16#0D#),
      1461 => to_slv(opcode_type, 16#07#),
      1462 => to_slv(opcode_type, 16#0F#),
      1463 => to_slv(opcode_type, 16#0A#),
      1464 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#06#),
      1473 => to_slv(opcode_type, 16#02#),
      1474 => to_slv(opcode_type, 16#06#),
      1475 => to_slv(opcode_type, 16#07#),
      1476 => to_slv(opcode_type, 16#0E#),
      1477 => to_slv(opcode_type, 16#11#),
      1478 => to_slv(opcode_type, 16#06#),
      1479 => to_slv(opcode_type, 16#0E#),
      1480 => to_slv(opcode_type, 16#10#),
      1481 => to_slv(opcode_type, 16#06#),
      1482 => to_slv(opcode_type, 16#07#),
      1483 => to_slv(opcode_type, 16#07#),
      1484 => to_slv(opcode_type, 16#0C#),
      1485 => to_slv(opcode_type, 16#5A#),
      1486 => to_slv(opcode_type, 16#06#),
      1487 => to_slv(opcode_type, 16#0A#),
      1488 => to_slv(opcode_type, 16#0B#),
      1489 => to_slv(opcode_type, 16#07#),
      1490 => to_slv(opcode_type, 16#09#),
      1491 => to_slv(opcode_type, 16#0F#),
      1492 => to_slv(opcode_type, 16#0C#),
      1493 => to_slv(opcode_type, 16#07#),
      1494 => to_slv(opcode_type, 16#0E#),
      1495 => to_slv(opcode_type, 16#0D#),
      1496 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#06#),
      1505 => to_slv(opcode_type, 16#03#),
      1506 => to_slv(opcode_type, 16#09#),
      1507 => to_slv(opcode_type, 16#07#),
      1508 => to_slv(opcode_type, 16#0D#),
      1509 => to_slv(opcode_type, 16#0E#),
      1510 => to_slv(opcode_type, 16#08#),
      1511 => to_slv(opcode_type, 16#10#),
      1512 => to_slv(opcode_type, 16#11#),
      1513 => to_slv(opcode_type, 16#06#),
      1514 => to_slv(opcode_type, 16#07#),
      1515 => to_slv(opcode_type, 16#07#),
      1516 => to_slv(opcode_type, 16#0B#),
      1517 => to_slv(opcode_type, 16#10#),
      1518 => to_slv(opcode_type, 16#07#),
      1519 => to_slv(opcode_type, 16#0A#),
      1520 => to_slv(opcode_type, 16#0E#),
      1521 => to_slv(opcode_type, 16#07#),
      1522 => to_slv(opcode_type, 16#07#),
      1523 => to_slv(opcode_type, 16#0A#),
      1524 => to_slv(opcode_type, 16#0B#),
      1525 => to_slv(opcode_type, 16#09#),
      1526 => to_slv(opcode_type, 16#59#),
      1527 => to_slv(opcode_type, 16#D8#),
      1528 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#07#),
      1537 => to_slv(opcode_type, 16#04#),
      1538 => to_slv(opcode_type, 16#06#),
      1539 => to_slv(opcode_type, 16#07#),
      1540 => to_slv(opcode_type, 16#11#),
      1541 => to_slv(opcode_type, 16#11#),
      1542 => to_slv(opcode_type, 16#09#),
      1543 => to_slv(opcode_type, 16#0E#),
      1544 => to_slv(opcode_type, 16#0E#),
      1545 => to_slv(opcode_type, 16#09#),
      1546 => to_slv(opcode_type, 16#08#),
      1547 => to_slv(opcode_type, 16#06#),
      1548 => to_slv(opcode_type, 16#0D#),
      1549 => to_slv(opcode_type, 16#0F#),
      1550 => to_slv(opcode_type, 16#08#),
      1551 => to_slv(opcode_type, 16#11#),
      1552 => to_slv(opcode_type, 16#A0#),
      1553 => to_slv(opcode_type, 16#08#),
      1554 => to_slv(opcode_type, 16#06#),
      1555 => to_slv(opcode_type, 16#2E#),
      1556 => to_slv(opcode_type, 16#0D#),
      1557 => to_slv(opcode_type, 16#08#),
      1558 => to_slv(opcode_type, 16#0C#),
      1559 => to_slv(opcode_type, 16#0E#),
      1560 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#08#),
      1569 => to_slv(opcode_type, 16#04#),
      1570 => to_slv(opcode_type, 16#09#),
      1571 => to_slv(opcode_type, 16#08#),
      1572 => to_slv(opcode_type, 16#0D#),
      1573 => to_slv(opcode_type, 16#0C#),
      1574 => to_slv(opcode_type, 16#07#),
      1575 => to_slv(opcode_type, 16#0F#),
      1576 => to_slv(opcode_type, 16#11#),
      1577 => to_slv(opcode_type, 16#09#),
      1578 => to_slv(opcode_type, 16#06#),
      1579 => to_slv(opcode_type, 16#07#),
      1580 => to_slv(opcode_type, 16#0F#),
      1581 => to_slv(opcode_type, 16#CF#),
      1582 => to_slv(opcode_type, 16#08#),
      1583 => to_slv(opcode_type, 16#0E#),
      1584 => to_slv(opcode_type, 16#0F#),
      1585 => to_slv(opcode_type, 16#08#),
      1586 => to_slv(opcode_type, 16#06#),
      1587 => to_slv(opcode_type, 16#0F#),
      1588 => to_slv(opcode_type, 16#11#),
      1589 => to_slv(opcode_type, 16#06#),
      1590 => to_slv(opcode_type, 16#0E#),
      1591 => to_slv(opcode_type, 16#10#),
      1592 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#08#),
      1601 => to_slv(opcode_type, 16#07#),
      1602 => to_slv(opcode_type, 16#04#),
      1603 => to_slv(opcode_type, 16#05#),
      1604 => to_slv(opcode_type, 16#0E#),
      1605 => to_slv(opcode_type, 16#09#),
      1606 => to_slv(opcode_type, 16#07#),
      1607 => to_slv(opcode_type, 16#10#),
      1608 => to_slv(opcode_type, 16#0B#),
      1609 => to_slv(opcode_type, 16#06#),
      1610 => to_slv(opcode_type, 16#10#),
      1611 => to_slv(opcode_type, 16#11#),
      1612 => to_slv(opcode_type, 16#06#),
      1613 => to_slv(opcode_type, 16#03#),
      1614 => to_slv(opcode_type, 16#06#),
      1615 => to_slv(opcode_type, 16#0A#),
      1616 => to_slv(opcode_type, 16#10#),
      1617 => to_slv(opcode_type, 16#09#),
      1618 => to_slv(opcode_type, 16#07#),
      1619 => to_slv(opcode_type, 16#0E#),
      1620 => to_slv(opcode_type, 16#0F#),
      1621 => to_slv(opcode_type, 16#06#),
      1622 => to_slv(opcode_type, 16#0D#),
      1623 => to_slv(opcode_type, 16#11#),
      1624 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#09#),
      1633 => to_slv(opcode_type, 16#06#),
      1634 => to_slv(opcode_type, 16#06#),
      1635 => to_slv(opcode_type, 16#07#),
      1636 => to_slv(opcode_type, 16#0E#),
      1637 => to_slv(opcode_type, 16#0D#),
      1638 => to_slv(opcode_type, 16#09#),
      1639 => to_slv(opcode_type, 16#0D#),
      1640 => to_slv(opcode_type, 16#0D#),
      1641 => to_slv(opcode_type, 16#06#),
      1642 => to_slv(opcode_type, 16#01#),
      1643 => to_slv(opcode_type, 16#0F#),
      1644 => to_slv(opcode_type, 16#01#),
      1645 => to_slv(opcode_type, 16#0E#),
      1646 => to_slv(opcode_type, 16#07#),
      1647 => to_slv(opcode_type, 16#02#),
      1648 => to_slv(opcode_type, 16#05#),
      1649 => to_slv(opcode_type, 16#11#),
      1650 => to_slv(opcode_type, 16#07#),
      1651 => to_slv(opcode_type, 16#01#),
      1652 => to_slv(opcode_type, 16#0B#),
      1653 => to_slv(opcode_type, 16#06#),
      1654 => to_slv(opcode_type, 16#0C#),
      1655 => to_slv(opcode_type, 16#0E#),
      1656 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#02#),
      1666 => to_slv(opcode_type, 16#06#),
      1667 => to_slv(opcode_type, 16#06#),
      1668 => to_slv(opcode_type, 16#10#),
      1669 => to_slv(opcode_type, 16#A8#),
      1670 => to_slv(opcode_type, 16#09#),
      1671 => to_slv(opcode_type, 16#0C#),
      1672 => to_slv(opcode_type, 16#0C#),
      1673 => to_slv(opcode_type, 16#09#),
      1674 => to_slv(opcode_type, 16#09#),
      1675 => to_slv(opcode_type, 16#09#),
      1676 => to_slv(opcode_type, 16#54#),
      1677 => to_slv(opcode_type, 16#10#),
      1678 => to_slv(opcode_type, 16#08#),
      1679 => to_slv(opcode_type, 16#0A#),
      1680 => to_slv(opcode_type, 16#10#),
      1681 => to_slv(opcode_type, 16#09#),
      1682 => to_slv(opcode_type, 16#06#),
      1683 => to_slv(opcode_type, 16#0D#),
      1684 => to_slv(opcode_type, 16#0E#),
      1685 => to_slv(opcode_type, 16#06#),
      1686 => to_slv(opcode_type, 16#F5#),
      1687 => to_slv(opcode_type, 16#0F#),
      1688 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#06#),
      1697 => to_slv(opcode_type, 16#02#),
      1698 => to_slv(opcode_type, 16#08#),
      1699 => to_slv(opcode_type, 16#09#),
      1700 => to_slv(opcode_type, 16#0F#),
      1701 => to_slv(opcode_type, 16#72#),
      1702 => to_slv(opcode_type, 16#07#),
      1703 => to_slv(opcode_type, 16#0C#),
      1704 => to_slv(opcode_type, 16#0B#),
      1705 => to_slv(opcode_type, 16#08#),
      1706 => to_slv(opcode_type, 16#09#),
      1707 => to_slv(opcode_type, 16#08#),
      1708 => to_slv(opcode_type, 16#0C#),
      1709 => to_slv(opcode_type, 16#92#),
      1710 => to_slv(opcode_type, 16#06#),
      1711 => to_slv(opcode_type, 16#0A#),
      1712 => to_slv(opcode_type, 16#0C#),
      1713 => to_slv(opcode_type, 16#06#),
      1714 => to_slv(opcode_type, 16#07#),
      1715 => to_slv(opcode_type, 16#10#),
      1716 => to_slv(opcode_type, 16#10#),
      1717 => to_slv(opcode_type, 16#07#),
      1718 => to_slv(opcode_type, 16#0B#),
      1719 => to_slv(opcode_type, 16#0C#),
      1720 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#09#),
      1729 => to_slv(opcode_type, 16#04#),
      1730 => to_slv(opcode_type, 16#07#),
      1731 => to_slv(opcode_type, 16#09#),
      1732 => to_slv(opcode_type, 16#58#),
      1733 => to_slv(opcode_type, 16#0D#),
      1734 => to_slv(opcode_type, 16#07#),
      1735 => to_slv(opcode_type, 16#0F#),
      1736 => to_slv(opcode_type, 16#11#),
      1737 => to_slv(opcode_type, 16#08#),
      1738 => to_slv(opcode_type, 16#06#),
      1739 => to_slv(opcode_type, 16#06#),
      1740 => to_slv(opcode_type, 16#0B#),
      1741 => to_slv(opcode_type, 16#11#),
      1742 => to_slv(opcode_type, 16#06#),
      1743 => to_slv(opcode_type, 16#0B#),
      1744 => to_slv(opcode_type, 16#0B#),
      1745 => to_slv(opcode_type, 16#08#),
      1746 => to_slv(opcode_type, 16#06#),
      1747 => to_slv(opcode_type, 16#11#),
      1748 => to_slv(opcode_type, 16#11#),
      1749 => to_slv(opcode_type, 16#07#),
      1750 => to_slv(opcode_type, 16#0D#),
      1751 => to_slv(opcode_type, 16#0F#),
      1752 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#09#),
      1761 => to_slv(opcode_type, 16#04#),
      1762 => to_slv(opcode_type, 16#09#),
      1763 => to_slv(opcode_type, 16#09#),
      1764 => to_slv(opcode_type, 16#10#),
      1765 => to_slv(opcode_type, 16#0F#),
      1766 => to_slv(opcode_type, 16#06#),
      1767 => to_slv(opcode_type, 16#1D#),
      1768 => to_slv(opcode_type, 16#0C#),
      1769 => to_slv(opcode_type, 16#08#),
      1770 => to_slv(opcode_type, 16#08#),
      1771 => to_slv(opcode_type, 16#07#),
      1772 => to_slv(opcode_type, 16#0B#),
      1773 => to_slv(opcode_type, 16#0E#),
      1774 => to_slv(opcode_type, 16#08#),
      1775 => to_slv(opcode_type, 16#0D#),
      1776 => to_slv(opcode_type, 16#0D#),
      1777 => to_slv(opcode_type, 16#09#),
      1778 => to_slv(opcode_type, 16#08#),
      1779 => to_slv(opcode_type, 16#0A#),
      1780 => to_slv(opcode_type, 16#0B#),
      1781 => to_slv(opcode_type, 16#09#),
      1782 => to_slv(opcode_type, 16#0D#),
      1783 => to_slv(opcode_type, 16#44#),
      1784 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#08#),
      1793 => to_slv(opcode_type, 16#03#),
      1794 => to_slv(opcode_type, 16#07#),
      1795 => to_slv(opcode_type, 16#07#),
      1796 => to_slv(opcode_type, 16#10#),
      1797 => to_slv(opcode_type, 16#0E#),
      1798 => to_slv(opcode_type, 16#06#),
      1799 => to_slv(opcode_type, 16#0C#),
      1800 => to_slv(opcode_type, 16#4C#),
      1801 => to_slv(opcode_type, 16#08#),
      1802 => to_slv(opcode_type, 16#06#),
      1803 => to_slv(opcode_type, 16#08#),
      1804 => to_slv(opcode_type, 16#0B#),
      1805 => to_slv(opcode_type, 16#0E#),
      1806 => to_slv(opcode_type, 16#09#),
      1807 => to_slv(opcode_type, 16#11#),
      1808 => to_slv(opcode_type, 16#0C#),
      1809 => to_slv(opcode_type, 16#07#),
      1810 => to_slv(opcode_type, 16#06#),
      1811 => to_slv(opcode_type, 16#11#),
      1812 => to_slv(opcode_type, 16#0E#),
      1813 => to_slv(opcode_type, 16#07#),
      1814 => to_slv(opcode_type, 16#0B#),
      1815 => to_slv(opcode_type, 16#10#),
      1816 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#08#),
      1825 => to_slv(opcode_type, 16#08#),
      1826 => to_slv(opcode_type, 16#05#),
      1827 => to_slv(opcode_type, 16#07#),
      1828 => to_slv(opcode_type, 16#11#),
      1829 => to_slv(opcode_type, 16#B5#),
      1830 => to_slv(opcode_type, 16#03#),
      1831 => to_slv(opcode_type, 16#01#),
      1832 => to_slv(opcode_type, 16#0F#),
      1833 => to_slv(opcode_type, 16#07#),
      1834 => to_slv(opcode_type, 16#06#),
      1835 => to_slv(opcode_type, 16#09#),
      1836 => to_slv(opcode_type, 16#0C#),
      1837 => to_slv(opcode_type, 16#0D#),
      1838 => to_slv(opcode_type, 16#08#),
      1839 => to_slv(opcode_type, 16#0F#),
      1840 => to_slv(opcode_type, 16#0F#),
      1841 => to_slv(opcode_type, 16#08#),
      1842 => to_slv(opcode_type, 16#08#),
      1843 => to_slv(opcode_type, 16#10#),
      1844 => to_slv(opcode_type, 16#D9#),
      1845 => to_slv(opcode_type, 16#09#),
      1846 => to_slv(opcode_type, 16#0A#),
      1847 => to_slv(opcode_type, 16#10#),
      1848 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#09#),
      1857 => to_slv(opcode_type, 16#04#),
      1858 => to_slv(opcode_type, 16#09#),
      1859 => to_slv(opcode_type, 16#07#),
      1860 => to_slv(opcode_type, 16#0C#),
      1861 => to_slv(opcode_type, 16#0F#),
      1862 => to_slv(opcode_type, 16#09#),
      1863 => to_slv(opcode_type, 16#0B#),
      1864 => to_slv(opcode_type, 16#0D#),
      1865 => to_slv(opcode_type, 16#09#),
      1866 => to_slv(opcode_type, 16#09#),
      1867 => to_slv(opcode_type, 16#06#),
      1868 => to_slv(opcode_type, 16#0D#),
      1869 => to_slv(opcode_type, 16#0B#),
      1870 => to_slv(opcode_type, 16#06#),
      1871 => to_slv(opcode_type, 16#8F#),
      1872 => to_slv(opcode_type, 16#41#),
      1873 => to_slv(opcode_type, 16#09#),
      1874 => to_slv(opcode_type, 16#08#),
      1875 => to_slv(opcode_type, 16#F9#),
      1876 => to_slv(opcode_type, 16#10#),
      1877 => to_slv(opcode_type, 16#08#),
      1878 => to_slv(opcode_type, 16#0A#),
      1879 => to_slv(opcode_type, 16#0E#),
      1880 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#08#),
      1889 => to_slv(opcode_type, 16#07#),
      1890 => to_slv(opcode_type, 16#02#),
      1891 => to_slv(opcode_type, 16#07#),
      1892 => to_slv(opcode_type, 16#0B#),
      1893 => to_slv(opcode_type, 16#35#),
      1894 => to_slv(opcode_type, 16#02#),
      1895 => to_slv(opcode_type, 16#01#),
      1896 => to_slv(opcode_type, 16#0E#),
      1897 => to_slv(opcode_type, 16#09#),
      1898 => to_slv(opcode_type, 16#08#),
      1899 => to_slv(opcode_type, 16#06#),
      1900 => to_slv(opcode_type, 16#0A#),
      1901 => to_slv(opcode_type, 16#0D#),
      1902 => to_slv(opcode_type, 16#08#),
      1903 => to_slv(opcode_type, 16#0C#),
      1904 => to_slv(opcode_type, 16#0C#),
      1905 => to_slv(opcode_type, 16#08#),
      1906 => to_slv(opcode_type, 16#08#),
      1907 => to_slv(opcode_type, 16#0A#),
      1908 => to_slv(opcode_type, 16#0A#),
      1909 => to_slv(opcode_type, 16#08#),
      1910 => to_slv(opcode_type, 16#0F#),
      1911 => to_slv(opcode_type, 16#D7#),
      1912 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#07#),
      1921 => to_slv(opcode_type, 16#09#),
      1922 => to_slv(opcode_type, 16#04#),
      1923 => to_slv(opcode_type, 16#05#),
      1924 => to_slv(opcode_type, 16#6E#),
      1925 => to_slv(opcode_type, 16#05#),
      1926 => to_slv(opcode_type, 16#07#),
      1927 => to_slv(opcode_type, 16#0C#),
      1928 => to_slv(opcode_type, 16#0B#),
      1929 => to_slv(opcode_type, 16#08#),
      1930 => to_slv(opcode_type, 16#06#),
      1931 => to_slv(opcode_type, 16#06#),
      1932 => to_slv(opcode_type, 16#0B#),
      1933 => to_slv(opcode_type, 16#0A#),
      1934 => to_slv(opcode_type, 16#07#),
      1935 => to_slv(opcode_type, 16#0F#),
      1936 => to_slv(opcode_type, 16#0B#),
      1937 => to_slv(opcode_type, 16#07#),
      1938 => to_slv(opcode_type, 16#09#),
      1939 => to_slv(opcode_type, 16#0B#),
      1940 => to_slv(opcode_type, 16#10#),
      1941 => to_slv(opcode_type, 16#09#),
      1942 => to_slv(opcode_type, 16#11#),
      1943 => to_slv(opcode_type, 16#0C#),
      1944 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#08#),
      1953 => to_slv(opcode_type, 16#06#),
      1954 => to_slv(opcode_type, 16#07#),
      1955 => to_slv(opcode_type, 16#04#),
      1956 => to_slv(opcode_type, 16#0E#),
      1957 => to_slv(opcode_type, 16#04#),
      1958 => to_slv(opcode_type, 16#11#),
      1959 => to_slv(opcode_type, 16#01#),
      1960 => to_slv(opcode_type, 16#07#),
      1961 => to_slv(opcode_type, 16#9B#),
      1962 => to_slv(opcode_type, 16#0C#),
      1963 => to_slv(opcode_type, 16#06#),
      1964 => to_slv(opcode_type, 16#06#),
      1965 => to_slv(opcode_type, 16#01#),
      1966 => to_slv(opcode_type, 16#11#),
      1967 => to_slv(opcode_type, 16#03#),
      1968 => to_slv(opcode_type, 16#0C#),
      1969 => to_slv(opcode_type, 16#08#),
      1970 => to_slv(opcode_type, 16#06#),
      1971 => to_slv(opcode_type, 16#0A#),
      1972 => to_slv(opcode_type, 16#10#),
      1973 => to_slv(opcode_type, 16#06#),
      1974 => to_slv(opcode_type, 16#0D#),
      1975 => to_slv(opcode_type, 16#0E#),
      1976 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#07#),
      1985 => to_slv(opcode_type, 16#01#),
      1986 => to_slv(opcode_type, 16#06#),
      1987 => to_slv(opcode_type, 16#09#),
      1988 => to_slv(opcode_type, 16#0B#),
      1989 => to_slv(opcode_type, 16#0A#),
      1990 => to_slv(opcode_type, 16#08#),
      1991 => to_slv(opcode_type, 16#0D#),
      1992 => to_slv(opcode_type, 16#11#),
      1993 => to_slv(opcode_type, 16#08#),
      1994 => to_slv(opcode_type, 16#08#),
      1995 => to_slv(opcode_type, 16#09#),
      1996 => to_slv(opcode_type, 16#10#),
      1997 => to_slv(opcode_type, 16#0C#),
      1998 => to_slv(opcode_type, 16#07#),
      1999 => to_slv(opcode_type, 16#10#),
      2000 => to_slv(opcode_type, 16#0B#),
      2001 => to_slv(opcode_type, 16#07#),
      2002 => to_slv(opcode_type, 16#09#),
      2003 => to_slv(opcode_type, 16#10#),
      2004 => to_slv(opcode_type, 16#0E#),
      2005 => to_slv(opcode_type, 16#08#),
      2006 => to_slv(opcode_type, 16#10#),
      2007 => to_slv(opcode_type, 16#11#),
      2008 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#07#),
      2017 => to_slv(opcode_type, 16#09#),
      2018 => to_slv(opcode_type, 16#03#),
      2019 => to_slv(opcode_type, 16#09#),
      2020 => to_slv(opcode_type, 16#0D#),
      2021 => to_slv(opcode_type, 16#0B#),
      2022 => to_slv(opcode_type, 16#08#),
      2023 => to_slv(opcode_type, 16#02#),
      2024 => to_slv(opcode_type, 16#0B#),
      2025 => to_slv(opcode_type, 16#06#),
      2026 => to_slv(opcode_type, 16#11#),
      2027 => to_slv(opcode_type, 16#0D#),
      2028 => to_slv(opcode_type, 16#07#),
      2029 => to_slv(opcode_type, 16#06#),
      2030 => to_slv(opcode_type, 16#09#),
      2031 => to_slv(opcode_type, 16#0E#),
      2032 => to_slv(opcode_type, 16#0A#),
      2033 => to_slv(opcode_type, 16#06#),
      2034 => to_slv(opcode_type, 16#61#),
      2035 => to_slv(opcode_type, 16#0A#),
      2036 => to_slv(opcode_type, 16#09#),
      2037 => to_slv(opcode_type, 16#03#),
      2038 => to_slv(opcode_type, 16#2E#),
      2039 => to_slv(opcode_type, 16#11#),
      2040 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#09#),
      2049 => to_slv(opcode_type, 16#01#),
      2050 => to_slv(opcode_type, 16#06#),
      2051 => to_slv(opcode_type, 16#07#),
      2052 => to_slv(opcode_type, 16#0D#),
      2053 => to_slv(opcode_type, 16#C5#),
      2054 => to_slv(opcode_type, 16#08#),
      2055 => to_slv(opcode_type, 16#10#),
      2056 => to_slv(opcode_type, 16#10#),
      2057 => to_slv(opcode_type, 16#08#),
      2058 => to_slv(opcode_type, 16#08#),
      2059 => to_slv(opcode_type, 16#07#),
      2060 => to_slv(opcode_type, 16#0E#),
      2061 => to_slv(opcode_type, 16#0E#),
      2062 => to_slv(opcode_type, 16#06#),
      2063 => to_slv(opcode_type, 16#0E#),
      2064 => to_slv(opcode_type, 16#10#),
      2065 => to_slv(opcode_type, 16#09#),
      2066 => to_slv(opcode_type, 16#06#),
      2067 => to_slv(opcode_type, 16#0D#),
      2068 => to_slv(opcode_type, 16#0C#),
      2069 => to_slv(opcode_type, 16#09#),
      2070 => to_slv(opcode_type, 16#0F#),
      2071 => to_slv(opcode_type, 16#0D#),
      2072 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#08#),
      2081 => to_slv(opcode_type, 16#03#),
      2082 => to_slv(opcode_type, 16#08#),
      2083 => to_slv(opcode_type, 16#09#),
      2084 => to_slv(opcode_type, 16#10#),
      2085 => to_slv(opcode_type, 16#0B#),
      2086 => to_slv(opcode_type, 16#08#),
      2087 => to_slv(opcode_type, 16#48#),
      2088 => to_slv(opcode_type, 16#0B#),
      2089 => to_slv(opcode_type, 16#07#),
      2090 => to_slv(opcode_type, 16#08#),
      2091 => to_slv(opcode_type, 16#08#),
      2092 => to_slv(opcode_type, 16#0C#),
      2093 => to_slv(opcode_type, 16#11#),
      2094 => to_slv(opcode_type, 16#06#),
      2095 => to_slv(opcode_type, 16#11#),
      2096 => to_slv(opcode_type, 16#11#),
      2097 => to_slv(opcode_type, 16#06#),
      2098 => to_slv(opcode_type, 16#09#),
      2099 => to_slv(opcode_type, 16#11#),
      2100 => to_slv(opcode_type, 16#0D#),
      2101 => to_slv(opcode_type, 16#07#),
      2102 => to_slv(opcode_type, 16#0F#),
      2103 => to_slv(opcode_type, 16#0C#),
      2104 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#07#),
      2113 => to_slv(opcode_type, 16#07#),
      2114 => to_slv(opcode_type, 16#05#),
      2115 => to_slv(opcode_type, 16#08#),
      2116 => to_slv(opcode_type, 16#0D#),
      2117 => to_slv(opcode_type, 16#0D#),
      2118 => to_slv(opcode_type, 16#07#),
      2119 => to_slv(opcode_type, 16#02#),
      2120 => to_slv(opcode_type, 16#0E#),
      2121 => to_slv(opcode_type, 16#06#),
      2122 => to_slv(opcode_type, 16#0B#),
      2123 => to_slv(opcode_type, 16#0D#),
      2124 => to_slv(opcode_type, 16#06#),
      2125 => to_slv(opcode_type, 16#07#),
      2126 => to_slv(opcode_type, 16#07#),
      2127 => to_slv(opcode_type, 16#0B#),
      2128 => to_slv(opcode_type, 16#0F#),
      2129 => to_slv(opcode_type, 16#02#),
      2130 => to_slv(opcode_type, 16#0D#),
      2131 => to_slv(opcode_type, 16#07#),
      2132 => to_slv(opcode_type, 16#01#),
      2133 => to_slv(opcode_type, 16#0A#),
      2134 => to_slv(opcode_type, 16#02#),
      2135 => to_slv(opcode_type, 16#10#),
      2136 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#08#),
      2145 => to_slv(opcode_type, 16#02#),
      2146 => to_slv(opcode_type, 16#09#),
      2147 => to_slv(opcode_type, 16#08#),
      2148 => to_slv(opcode_type, 16#0E#),
      2149 => to_slv(opcode_type, 16#10#),
      2150 => to_slv(opcode_type, 16#08#),
      2151 => to_slv(opcode_type, 16#0B#),
      2152 => to_slv(opcode_type, 16#0E#),
      2153 => to_slv(opcode_type, 16#09#),
      2154 => to_slv(opcode_type, 16#08#),
      2155 => to_slv(opcode_type, 16#08#),
      2156 => to_slv(opcode_type, 16#0A#),
      2157 => to_slv(opcode_type, 16#0D#),
      2158 => to_slv(opcode_type, 16#09#),
      2159 => to_slv(opcode_type, 16#11#),
      2160 => to_slv(opcode_type, 16#0B#),
      2161 => to_slv(opcode_type, 16#08#),
      2162 => to_slv(opcode_type, 16#08#),
      2163 => to_slv(opcode_type, 16#FA#),
      2164 => to_slv(opcode_type, 16#0E#),
      2165 => to_slv(opcode_type, 16#06#),
      2166 => to_slv(opcode_type, 16#0C#),
      2167 => to_slv(opcode_type, 16#11#),
      2168 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#07#),
      2177 => to_slv(opcode_type, 16#07#),
      2178 => to_slv(opcode_type, 16#04#),
      2179 => to_slv(opcode_type, 16#09#),
      2180 => to_slv(opcode_type, 16#10#),
      2181 => to_slv(opcode_type, 16#FC#),
      2182 => to_slv(opcode_type, 16#08#),
      2183 => to_slv(opcode_type, 16#09#),
      2184 => to_slv(opcode_type, 16#10#),
      2185 => to_slv(opcode_type, 16#11#),
      2186 => to_slv(opcode_type, 16#02#),
      2187 => to_slv(opcode_type, 16#0C#),
      2188 => to_slv(opcode_type, 16#06#),
      2189 => to_slv(opcode_type, 16#02#),
      2190 => to_slv(opcode_type, 16#07#),
      2191 => to_slv(opcode_type, 16#0B#),
      2192 => to_slv(opcode_type, 16#0C#),
      2193 => to_slv(opcode_type, 16#09#),
      2194 => to_slv(opcode_type, 16#09#),
      2195 => to_slv(opcode_type, 16#11#),
      2196 => to_slv(opcode_type, 16#10#),
      2197 => to_slv(opcode_type, 16#07#),
      2198 => to_slv(opcode_type, 16#0F#),
      2199 => to_slv(opcode_type, 16#11#),
      2200 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#09#),
      2209 => to_slv(opcode_type, 16#05#),
      2210 => to_slv(opcode_type, 16#06#),
      2211 => to_slv(opcode_type, 16#09#),
      2212 => to_slv(opcode_type, 16#10#),
      2213 => to_slv(opcode_type, 16#10#),
      2214 => to_slv(opcode_type, 16#06#),
      2215 => to_slv(opcode_type, 16#0E#),
      2216 => to_slv(opcode_type, 16#0A#),
      2217 => to_slv(opcode_type, 16#09#),
      2218 => to_slv(opcode_type, 16#07#),
      2219 => to_slv(opcode_type, 16#08#),
      2220 => to_slv(opcode_type, 16#0D#),
      2221 => to_slv(opcode_type, 16#0B#),
      2222 => to_slv(opcode_type, 16#07#),
      2223 => to_slv(opcode_type, 16#0E#),
      2224 => to_slv(opcode_type, 16#0B#),
      2225 => to_slv(opcode_type, 16#06#),
      2226 => to_slv(opcode_type, 16#06#),
      2227 => to_slv(opcode_type, 16#0A#),
      2228 => to_slv(opcode_type, 16#25#),
      2229 => to_slv(opcode_type, 16#06#),
      2230 => to_slv(opcode_type, 16#0E#),
      2231 => to_slv(opcode_type, 16#0E#),
      2232 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#05#),
      2242 => to_slv(opcode_type, 16#09#),
      2243 => to_slv(opcode_type, 16#08#),
      2244 => to_slv(opcode_type, 16#3C#),
      2245 => to_slv(opcode_type, 16#69#),
      2246 => to_slv(opcode_type, 16#06#),
      2247 => to_slv(opcode_type, 16#10#),
      2248 => to_slv(opcode_type, 16#0F#),
      2249 => to_slv(opcode_type, 16#07#),
      2250 => to_slv(opcode_type, 16#07#),
      2251 => to_slv(opcode_type, 16#08#),
      2252 => to_slv(opcode_type, 16#0C#),
      2253 => to_slv(opcode_type, 16#0D#),
      2254 => to_slv(opcode_type, 16#08#),
      2255 => to_slv(opcode_type, 16#0A#),
      2256 => to_slv(opcode_type, 16#0A#),
      2257 => to_slv(opcode_type, 16#09#),
      2258 => to_slv(opcode_type, 16#08#),
      2259 => to_slv(opcode_type, 16#0F#),
      2260 => to_slv(opcode_type, 16#0C#),
      2261 => to_slv(opcode_type, 16#09#),
      2262 => to_slv(opcode_type, 16#10#),
      2263 => to_slv(opcode_type, 16#10#),
      2264 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#07#),
      2273 => to_slv(opcode_type, 16#07#),
      2274 => to_slv(opcode_type, 16#07#),
      2275 => to_slv(opcode_type, 16#01#),
      2276 => to_slv(opcode_type, 16#0F#),
      2277 => to_slv(opcode_type, 16#03#),
      2278 => to_slv(opcode_type, 16#0C#),
      2279 => to_slv(opcode_type, 16#08#),
      2280 => to_slv(opcode_type, 16#05#),
      2281 => to_slv(opcode_type, 16#0E#),
      2282 => to_slv(opcode_type, 16#01#),
      2283 => to_slv(opcode_type, 16#0B#),
      2284 => to_slv(opcode_type, 16#09#),
      2285 => to_slv(opcode_type, 16#09#),
      2286 => to_slv(opcode_type, 16#02#),
      2287 => to_slv(opcode_type, 16#11#),
      2288 => to_slv(opcode_type, 16#08#),
      2289 => to_slv(opcode_type, 16#0A#),
      2290 => to_slv(opcode_type, 16#0E#),
      2291 => to_slv(opcode_type, 16#06#),
      2292 => to_slv(opcode_type, 16#07#),
      2293 => to_slv(opcode_type, 16#0D#),
      2294 => to_slv(opcode_type, 16#10#),
      2295 => to_slv(opcode_type, 16#11#),
      2296 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#06#),
      2305 => to_slv(opcode_type, 16#05#),
      2306 => to_slv(opcode_type, 16#06#),
      2307 => to_slv(opcode_type, 16#09#),
      2308 => to_slv(opcode_type, 16#0B#),
      2309 => to_slv(opcode_type, 16#0F#),
      2310 => to_slv(opcode_type, 16#06#),
      2311 => to_slv(opcode_type, 16#0B#),
      2312 => to_slv(opcode_type, 16#0A#),
      2313 => to_slv(opcode_type, 16#08#),
      2314 => to_slv(opcode_type, 16#08#),
      2315 => to_slv(opcode_type, 16#09#),
      2316 => to_slv(opcode_type, 16#11#),
      2317 => to_slv(opcode_type, 16#3B#),
      2318 => to_slv(opcode_type, 16#07#),
      2319 => to_slv(opcode_type, 16#0A#),
      2320 => to_slv(opcode_type, 16#11#),
      2321 => to_slv(opcode_type, 16#09#),
      2322 => to_slv(opcode_type, 16#07#),
      2323 => to_slv(opcode_type, 16#0C#),
      2324 => to_slv(opcode_type, 16#0A#),
      2325 => to_slv(opcode_type, 16#09#),
      2326 => to_slv(opcode_type, 16#0E#),
      2327 => to_slv(opcode_type, 16#0E#),
      2328 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#06#),
      2337 => to_slv(opcode_type, 16#02#),
      2338 => to_slv(opcode_type, 16#08#),
      2339 => to_slv(opcode_type, 16#07#),
      2340 => to_slv(opcode_type, 16#0C#),
      2341 => to_slv(opcode_type, 16#11#),
      2342 => to_slv(opcode_type, 16#09#),
      2343 => to_slv(opcode_type, 16#0D#),
      2344 => to_slv(opcode_type, 16#0C#),
      2345 => to_slv(opcode_type, 16#09#),
      2346 => to_slv(opcode_type, 16#09#),
      2347 => to_slv(opcode_type, 16#06#),
      2348 => to_slv(opcode_type, 16#0D#),
      2349 => to_slv(opcode_type, 16#0B#),
      2350 => to_slv(opcode_type, 16#08#),
      2351 => to_slv(opcode_type, 16#11#),
      2352 => to_slv(opcode_type, 16#AC#),
      2353 => to_slv(opcode_type, 16#09#),
      2354 => to_slv(opcode_type, 16#08#),
      2355 => to_slv(opcode_type, 16#0F#),
      2356 => to_slv(opcode_type, 16#10#),
      2357 => to_slv(opcode_type, 16#06#),
      2358 => to_slv(opcode_type, 16#0A#),
      2359 => to_slv(opcode_type, 16#0F#),
      2360 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#06#),
      2369 => to_slv(opcode_type, 16#07#),
      2370 => to_slv(opcode_type, 16#03#),
      2371 => to_slv(opcode_type, 16#07#),
      2372 => to_slv(opcode_type, 16#0B#),
      2373 => to_slv(opcode_type, 16#10#),
      2374 => to_slv(opcode_type, 16#02#),
      2375 => to_slv(opcode_type, 16#09#),
      2376 => to_slv(opcode_type, 16#10#),
      2377 => to_slv(opcode_type, 16#0D#),
      2378 => to_slv(opcode_type, 16#06#),
      2379 => to_slv(opcode_type, 16#07#),
      2380 => to_slv(opcode_type, 16#04#),
      2381 => to_slv(opcode_type, 16#11#),
      2382 => to_slv(opcode_type, 16#08#),
      2383 => to_slv(opcode_type, 16#0B#),
      2384 => to_slv(opcode_type, 16#0F#),
      2385 => to_slv(opcode_type, 16#08#),
      2386 => to_slv(opcode_type, 16#07#),
      2387 => to_slv(opcode_type, 16#11#),
      2388 => to_slv(opcode_type, 16#0C#),
      2389 => to_slv(opcode_type, 16#07#),
      2390 => to_slv(opcode_type, 16#11#),
      2391 => to_slv(opcode_type, 16#77#),
      2392 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#09#),
      2401 => to_slv(opcode_type, 16#09#),
      2402 => to_slv(opcode_type, 16#02#),
      2403 => to_slv(opcode_type, 16#07#),
      2404 => to_slv(opcode_type, 16#0F#),
      2405 => to_slv(opcode_type, 16#11#),
      2406 => to_slv(opcode_type, 16#07#),
      2407 => to_slv(opcode_type, 16#09#),
      2408 => to_slv(opcode_type, 16#93#),
      2409 => to_slv(opcode_type, 16#11#),
      2410 => to_slv(opcode_type, 16#04#),
      2411 => to_slv(opcode_type, 16#0C#),
      2412 => to_slv(opcode_type, 16#08#),
      2413 => to_slv(opcode_type, 16#02#),
      2414 => to_slv(opcode_type, 16#07#),
      2415 => to_slv(opcode_type, 16#0C#),
      2416 => to_slv(opcode_type, 16#0A#),
      2417 => to_slv(opcode_type, 16#09#),
      2418 => to_slv(opcode_type, 16#08#),
      2419 => to_slv(opcode_type, 16#0E#),
      2420 => to_slv(opcode_type, 16#10#),
      2421 => to_slv(opcode_type, 16#09#),
      2422 => to_slv(opcode_type, 16#0E#),
      2423 => to_slv(opcode_type, 16#0E#),
      2424 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#09#),
      2433 => to_slv(opcode_type, 16#08#),
      2434 => to_slv(opcode_type, 16#05#),
      2435 => to_slv(opcode_type, 16#05#),
      2436 => to_slv(opcode_type, 16#0F#),
      2437 => to_slv(opcode_type, 16#04#),
      2438 => to_slv(opcode_type, 16#08#),
      2439 => to_slv(opcode_type, 16#0F#),
      2440 => to_slv(opcode_type, 16#0E#),
      2441 => to_slv(opcode_type, 16#06#),
      2442 => to_slv(opcode_type, 16#08#),
      2443 => to_slv(opcode_type, 16#06#),
      2444 => to_slv(opcode_type, 16#0F#),
      2445 => to_slv(opcode_type, 16#AF#),
      2446 => to_slv(opcode_type, 16#07#),
      2447 => to_slv(opcode_type, 16#0B#),
      2448 => to_slv(opcode_type, 16#0A#),
      2449 => to_slv(opcode_type, 16#09#),
      2450 => to_slv(opcode_type, 16#09#),
      2451 => to_slv(opcode_type, 16#0C#),
      2452 => to_slv(opcode_type, 16#65#),
      2453 => to_slv(opcode_type, 16#09#),
      2454 => to_slv(opcode_type, 16#11#),
      2455 => to_slv(opcode_type, 16#10#),
      2456 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#09#),
      2465 => to_slv(opcode_type, 16#02#),
      2466 => to_slv(opcode_type, 16#09#),
      2467 => to_slv(opcode_type, 16#06#),
      2468 => to_slv(opcode_type, 16#0B#),
      2469 => to_slv(opcode_type, 16#0A#),
      2470 => to_slv(opcode_type, 16#06#),
      2471 => to_slv(opcode_type, 16#11#),
      2472 => to_slv(opcode_type, 16#0C#),
      2473 => to_slv(opcode_type, 16#07#),
      2474 => to_slv(opcode_type, 16#06#),
      2475 => to_slv(opcode_type, 16#06#),
      2476 => to_slv(opcode_type, 16#0E#),
      2477 => to_slv(opcode_type, 16#11#),
      2478 => to_slv(opcode_type, 16#06#),
      2479 => to_slv(opcode_type, 16#11#),
      2480 => to_slv(opcode_type, 16#0E#),
      2481 => to_slv(opcode_type, 16#06#),
      2482 => to_slv(opcode_type, 16#09#),
      2483 => to_slv(opcode_type, 16#0C#),
      2484 => to_slv(opcode_type, 16#10#),
      2485 => to_slv(opcode_type, 16#08#),
      2486 => to_slv(opcode_type, 16#0C#),
      2487 => to_slv(opcode_type, 16#0F#),
      2488 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#08#),
      2497 => to_slv(opcode_type, 16#02#),
      2498 => to_slv(opcode_type, 16#09#),
      2499 => to_slv(opcode_type, 16#06#),
      2500 => to_slv(opcode_type, 16#0D#),
      2501 => to_slv(opcode_type, 16#0A#),
      2502 => to_slv(opcode_type, 16#08#),
      2503 => to_slv(opcode_type, 16#9C#),
      2504 => to_slv(opcode_type, 16#0E#),
      2505 => to_slv(opcode_type, 16#07#),
      2506 => to_slv(opcode_type, 16#06#),
      2507 => to_slv(opcode_type, 16#07#),
      2508 => to_slv(opcode_type, 16#10#),
      2509 => to_slv(opcode_type, 16#0F#),
      2510 => to_slv(opcode_type, 16#06#),
      2511 => to_slv(opcode_type, 16#0B#),
      2512 => to_slv(opcode_type, 16#10#),
      2513 => to_slv(opcode_type, 16#09#),
      2514 => to_slv(opcode_type, 16#06#),
      2515 => to_slv(opcode_type, 16#0F#),
      2516 => to_slv(opcode_type, 16#0D#),
      2517 => to_slv(opcode_type, 16#06#),
      2518 => to_slv(opcode_type, 16#0A#),
      2519 => to_slv(opcode_type, 16#0A#),
      2520 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#09#),
      2529 => to_slv(opcode_type, 16#04#),
      2530 => to_slv(opcode_type, 16#06#),
      2531 => to_slv(opcode_type, 16#08#),
      2532 => to_slv(opcode_type, 16#0F#),
      2533 => to_slv(opcode_type, 16#0A#),
      2534 => to_slv(opcode_type, 16#09#),
      2535 => to_slv(opcode_type, 16#0B#),
      2536 => to_slv(opcode_type, 16#10#),
      2537 => to_slv(opcode_type, 16#07#),
      2538 => to_slv(opcode_type, 16#07#),
      2539 => to_slv(opcode_type, 16#06#),
      2540 => to_slv(opcode_type, 16#0E#),
      2541 => to_slv(opcode_type, 16#0D#),
      2542 => to_slv(opcode_type, 16#07#),
      2543 => to_slv(opcode_type, 16#0B#),
      2544 => to_slv(opcode_type, 16#0F#),
      2545 => to_slv(opcode_type, 16#06#),
      2546 => to_slv(opcode_type, 16#07#),
      2547 => to_slv(opcode_type, 16#0E#),
      2548 => to_slv(opcode_type, 16#0D#),
      2549 => to_slv(opcode_type, 16#08#),
      2550 => to_slv(opcode_type, 16#11#),
      2551 => to_slv(opcode_type, 16#1F#),
      2552 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#09#),
      2561 => to_slv(opcode_type, 16#02#),
      2562 => to_slv(opcode_type, 16#08#),
      2563 => to_slv(opcode_type, 16#06#),
      2564 => to_slv(opcode_type, 16#0A#),
      2565 => to_slv(opcode_type, 16#0C#),
      2566 => to_slv(opcode_type, 16#07#),
      2567 => to_slv(opcode_type, 16#10#),
      2568 => to_slv(opcode_type, 16#0A#),
      2569 => to_slv(opcode_type, 16#08#),
      2570 => to_slv(opcode_type, 16#09#),
      2571 => to_slv(opcode_type, 16#06#),
      2572 => to_slv(opcode_type, 16#11#),
      2573 => to_slv(opcode_type, 16#CC#),
      2574 => to_slv(opcode_type, 16#09#),
      2575 => to_slv(opcode_type, 16#0C#),
      2576 => to_slv(opcode_type, 16#0D#),
      2577 => to_slv(opcode_type, 16#07#),
      2578 => to_slv(opcode_type, 16#08#),
      2579 => to_slv(opcode_type, 16#0F#),
      2580 => to_slv(opcode_type, 16#11#),
      2581 => to_slv(opcode_type, 16#06#),
      2582 => to_slv(opcode_type, 16#0E#),
      2583 => to_slv(opcode_type, 16#0F#),
      2584 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#08#),
      2593 => to_slv(opcode_type, 16#08#),
      2594 => to_slv(opcode_type, 16#04#),
      2595 => to_slv(opcode_type, 16#02#),
      2596 => to_slv(opcode_type, 16#0A#),
      2597 => to_slv(opcode_type, 16#04#),
      2598 => to_slv(opcode_type, 16#06#),
      2599 => to_slv(opcode_type, 16#0F#),
      2600 => to_slv(opcode_type, 16#0C#),
      2601 => to_slv(opcode_type, 16#08#),
      2602 => to_slv(opcode_type, 16#09#),
      2603 => to_slv(opcode_type, 16#06#),
      2604 => to_slv(opcode_type, 16#0E#),
      2605 => to_slv(opcode_type, 16#0B#),
      2606 => to_slv(opcode_type, 16#06#),
      2607 => to_slv(opcode_type, 16#0E#),
      2608 => to_slv(opcode_type, 16#10#),
      2609 => to_slv(opcode_type, 16#07#),
      2610 => to_slv(opcode_type, 16#07#),
      2611 => to_slv(opcode_type, 16#0E#),
      2612 => to_slv(opcode_type, 16#0D#),
      2613 => to_slv(opcode_type, 16#07#),
      2614 => to_slv(opcode_type, 16#0D#),
      2615 => to_slv(opcode_type, 16#11#),
      2616 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#06#),
      2625 => to_slv(opcode_type, 16#05#),
      2626 => to_slv(opcode_type, 16#09#),
      2627 => to_slv(opcode_type, 16#09#),
      2628 => to_slv(opcode_type, 16#0A#),
      2629 => to_slv(opcode_type, 16#0C#),
      2630 => to_slv(opcode_type, 16#07#),
      2631 => to_slv(opcode_type, 16#0B#),
      2632 => to_slv(opcode_type, 16#0B#),
      2633 => to_slv(opcode_type, 16#07#),
      2634 => to_slv(opcode_type, 16#08#),
      2635 => to_slv(opcode_type, 16#07#),
      2636 => to_slv(opcode_type, 16#0D#),
      2637 => to_slv(opcode_type, 16#0A#),
      2638 => to_slv(opcode_type, 16#08#),
      2639 => to_slv(opcode_type, 16#0A#),
      2640 => to_slv(opcode_type, 16#0E#),
      2641 => to_slv(opcode_type, 16#08#),
      2642 => to_slv(opcode_type, 16#08#),
      2643 => to_slv(opcode_type, 16#10#),
      2644 => to_slv(opcode_type, 16#B6#),
      2645 => to_slv(opcode_type, 16#06#),
      2646 => to_slv(opcode_type, 16#0C#),
      2647 => to_slv(opcode_type, 16#0B#),
      2648 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#06#),
      2657 => to_slv(opcode_type, 16#08#),
      2658 => to_slv(opcode_type, 16#08#),
      2659 => to_slv(opcode_type, 16#09#),
      2660 => to_slv(opcode_type, 16#0A#),
      2661 => to_slv(opcode_type, 16#0E#),
      2662 => to_slv(opcode_type, 16#01#),
      2663 => to_slv(opcode_type, 16#0E#),
      2664 => to_slv(opcode_type, 16#01#),
      2665 => to_slv(opcode_type, 16#01#),
      2666 => to_slv(opcode_type, 16#0A#),
      2667 => to_slv(opcode_type, 16#09#),
      2668 => to_slv(opcode_type, 16#08#),
      2669 => to_slv(opcode_type, 16#03#),
      2670 => to_slv(opcode_type, 16#0F#),
      2671 => to_slv(opcode_type, 16#06#),
      2672 => to_slv(opcode_type, 16#0A#),
      2673 => to_slv(opcode_type, 16#0C#),
      2674 => to_slv(opcode_type, 16#08#),
      2675 => to_slv(opcode_type, 16#07#),
      2676 => to_slv(opcode_type, 16#0D#),
      2677 => to_slv(opcode_type, 16#10#),
      2678 => to_slv(opcode_type, 16#02#),
      2679 => to_slv(opcode_type, 16#0F#),
      2680 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#06#),
      2689 => to_slv(opcode_type, 16#05#),
      2690 => to_slv(opcode_type, 16#07#),
      2691 => to_slv(opcode_type, 16#08#),
      2692 => to_slv(opcode_type, 16#0B#),
      2693 => to_slv(opcode_type, 16#0D#),
      2694 => to_slv(opcode_type, 16#07#),
      2695 => to_slv(opcode_type, 16#0F#),
      2696 => to_slv(opcode_type, 16#0D#),
      2697 => to_slv(opcode_type, 16#08#),
      2698 => to_slv(opcode_type, 16#07#),
      2699 => to_slv(opcode_type, 16#08#),
      2700 => to_slv(opcode_type, 16#0A#),
      2701 => to_slv(opcode_type, 16#0B#),
      2702 => to_slv(opcode_type, 16#07#),
      2703 => to_slv(opcode_type, 16#0B#),
      2704 => to_slv(opcode_type, 16#94#),
      2705 => to_slv(opcode_type, 16#08#),
      2706 => to_slv(opcode_type, 16#08#),
      2707 => to_slv(opcode_type, 16#0C#),
      2708 => to_slv(opcode_type, 16#0B#),
      2709 => to_slv(opcode_type, 16#07#),
      2710 => to_slv(opcode_type, 16#10#),
      2711 => to_slv(opcode_type, 16#0B#),
      2712 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#08#),
      2721 => to_slv(opcode_type, 16#06#),
      2722 => to_slv(opcode_type, 16#04#),
      2723 => to_slv(opcode_type, 16#07#),
      2724 => to_slv(opcode_type, 16#0C#),
      2725 => to_slv(opcode_type, 16#84#),
      2726 => to_slv(opcode_type, 16#01#),
      2727 => to_slv(opcode_type, 16#08#),
      2728 => to_slv(opcode_type, 16#0D#),
      2729 => to_slv(opcode_type, 16#10#),
      2730 => to_slv(opcode_type, 16#06#),
      2731 => to_slv(opcode_type, 16#06#),
      2732 => to_slv(opcode_type, 16#04#),
      2733 => to_slv(opcode_type, 16#0F#),
      2734 => to_slv(opcode_type, 16#07#),
      2735 => to_slv(opcode_type, 16#0B#),
      2736 => to_slv(opcode_type, 16#0A#),
      2737 => to_slv(opcode_type, 16#09#),
      2738 => to_slv(opcode_type, 16#07#),
      2739 => to_slv(opcode_type, 16#0B#),
      2740 => to_slv(opcode_type, 16#72#),
      2741 => to_slv(opcode_type, 16#07#),
      2742 => to_slv(opcode_type, 16#0B#),
      2743 => to_slv(opcode_type, 16#0B#),
      2744 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#07#),
      2753 => to_slv(opcode_type, 16#01#),
      2754 => to_slv(opcode_type, 16#08#),
      2755 => to_slv(opcode_type, 16#09#),
      2756 => to_slv(opcode_type, 16#0F#),
      2757 => to_slv(opcode_type, 16#0B#),
      2758 => to_slv(opcode_type, 16#09#),
      2759 => to_slv(opcode_type, 16#0C#),
      2760 => to_slv(opcode_type, 16#0C#),
      2761 => to_slv(opcode_type, 16#09#),
      2762 => to_slv(opcode_type, 16#06#),
      2763 => to_slv(opcode_type, 16#07#),
      2764 => to_slv(opcode_type, 16#52#),
      2765 => to_slv(opcode_type, 16#10#),
      2766 => to_slv(opcode_type, 16#06#),
      2767 => to_slv(opcode_type, 16#11#),
      2768 => to_slv(opcode_type, 16#0C#),
      2769 => to_slv(opcode_type, 16#09#),
      2770 => to_slv(opcode_type, 16#06#),
      2771 => to_slv(opcode_type, 16#10#),
      2772 => to_slv(opcode_type, 16#0E#),
      2773 => to_slv(opcode_type, 16#06#),
      2774 => to_slv(opcode_type, 16#0B#),
      2775 => to_slv(opcode_type, 16#11#),
      2776 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#06#),
      2785 => to_slv(opcode_type, 16#02#),
      2786 => to_slv(opcode_type, 16#09#),
      2787 => to_slv(opcode_type, 16#06#),
      2788 => to_slv(opcode_type, 16#0F#),
      2789 => to_slv(opcode_type, 16#0B#),
      2790 => to_slv(opcode_type, 16#06#),
      2791 => to_slv(opcode_type, 16#0C#),
      2792 => to_slv(opcode_type, 16#0C#),
      2793 => to_slv(opcode_type, 16#07#),
      2794 => to_slv(opcode_type, 16#06#),
      2795 => to_slv(opcode_type, 16#07#),
      2796 => to_slv(opcode_type, 16#0F#),
      2797 => to_slv(opcode_type, 16#0A#),
      2798 => to_slv(opcode_type, 16#08#),
      2799 => to_slv(opcode_type, 16#B6#),
      2800 => to_slv(opcode_type, 16#0B#),
      2801 => to_slv(opcode_type, 16#09#),
      2802 => to_slv(opcode_type, 16#08#),
      2803 => to_slv(opcode_type, 16#10#),
      2804 => to_slv(opcode_type, 16#0F#),
      2805 => to_slv(opcode_type, 16#06#),
      2806 => to_slv(opcode_type, 16#79#),
      2807 => to_slv(opcode_type, 16#0A#),
      2808 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#09#),
      2817 => to_slv(opcode_type, 16#08#),
      2818 => to_slv(opcode_type, 16#01#),
      2819 => to_slv(opcode_type, 16#03#),
      2820 => to_slv(opcode_type, 16#0E#),
      2821 => to_slv(opcode_type, 16#06#),
      2822 => to_slv(opcode_type, 16#05#),
      2823 => to_slv(opcode_type, 16#0E#),
      2824 => to_slv(opcode_type, 16#03#),
      2825 => to_slv(opcode_type, 16#0A#),
      2826 => to_slv(opcode_type, 16#09#),
      2827 => to_slv(opcode_type, 16#09#),
      2828 => to_slv(opcode_type, 16#08#),
      2829 => to_slv(opcode_type, 16#0A#),
      2830 => to_slv(opcode_type, 16#0B#),
      2831 => to_slv(opcode_type, 16#05#),
      2832 => to_slv(opcode_type, 16#0A#),
      2833 => to_slv(opcode_type, 16#08#),
      2834 => to_slv(opcode_type, 16#09#),
      2835 => to_slv(opcode_type, 16#0B#),
      2836 => to_slv(opcode_type, 16#0B#),
      2837 => to_slv(opcode_type, 16#08#),
      2838 => to_slv(opcode_type, 16#0A#),
      2839 => to_slv(opcode_type, 16#0F#),
      2840 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#09#),
      2849 => to_slv(opcode_type, 16#05#),
      2850 => to_slv(opcode_type, 16#09#),
      2851 => to_slv(opcode_type, 16#09#),
      2852 => to_slv(opcode_type, 16#0E#),
      2853 => to_slv(opcode_type, 16#0E#),
      2854 => to_slv(opcode_type, 16#09#),
      2855 => to_slv(opcode_type, 16#5F#),
      2856 => to_slv(opcode_type, 16#DD#),
      2857 => to_slv(opcode_type, 16#08#),
      2858 => to_slv(opcode_type, 16#08#),
      2859 => to_slv(opcode_type, 16#07#),
      2860 => to_slv(opcode_type, 16#11#),
      2861 => to_slv(opcode_type, 16#0B#),
      2862 => to_slv(opcode_type, 16#08#),
      2863 => to_slv(opcode_type, 16#0F#),
      2864 => to_slv(opcode_type, 16#0A#),
      2865 => to_slv(opcode_type, 16#09#),
      2866 => to_slv(opcode_type, 16#09#),
      2867 => to_slv(opcode_type, 16#E9#),
      2868 => to_slv(opcode_type, 16#0A#),
      2869 => to_slv(opcode_type, 16#08#),
      2870 => to_slv(opcode_type, 16#10#),
      2871 => to_slv(opcode_type, 16#0B#),
      2872 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#08#),
      2881 => to_slv(opcode_type, 16#04#),
      2882 => to_slv(opcode_type, 16#07#),
      2883 => to_slv(opcode_type, 16#08#),
      2884 => to_slv(opcode_type, 16#0A#),
      2885 => to_slv(opcode_type, 16#0A#),
      2886 => to_slv(opcode_type, 16#07#),
      2887 => to_slv(opcode_type, 16#0A#),
      2888 => to_slv(opcode_type, 16#0B#),
      2889 => to_slv(opcode_type, 16#09#),
      2890 => to_slv(opcode_type, 16#06#),
      2891 => to_slv(opcode_type, 16#07#),
      2892 => to_slv(opcode_type, 16#50#),
      2893 => to_slv(opcode_type, 16#11#),
      2894 => to_slv(opcode_type, 16#09#),
      2895 => to_slv(opcode_type, 16#0D#),
      2896 => to_slv(opcode_type, 16#0D#),
      2897 => to_slv(opcode_type, 16#06#),
      2898 => to_slv(opcode_type, 16#09#),
      2899 => to_slv(opcode_type, 16#0C#),
      2900 => to_slv(opcode_type, 16#79#),
      2901 => to_slv(opcode_type, 16#09#),
      2902 => to_slv(opcode_type, 16#0F#),
      2903 => to_slv(opcode_type, 16#0F#),
      2904 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#06#),
      2913 => to_slv(opcode_type, 16#01#),
      2914 => to_slv(opcode_type, 16#08#),
      2915 => to_slv(opcode_type, 16#06#),
      2916 => to_slv(opcode_type, 16#E6#),
      2917 => to_slv(opcode_type, 16#9D#),
      2918 => to_slv(opcode_type, 16#09#),
      2919 => to_slv(opcode_type, 16#0B#),
      2920 => to_slv(opcode_type, 16#0A#),
      2921 => to_slv(opcode_type, 16#07#),
      2922 => to_slv(opcode_type, 16#09#),
      2923 => to_slv(opcode_type, 16#09#),
      2924 => to_slv(opcode_type, 16#0E#),
      2925 => to_slv(opcode_type, 16#0D#),
      2926 => to_slv(opcode_type, 16#08#),
      2927 => to_slv(opcode_type, 16#11#),
      2928 => to_slv(opcode_type, 16#10#),
      2929 => to_slv(opcode_type, 16#09#),
      2930 => to_slv(opcode_type, 16#06#),
      2931 => to_slv(opcode_type, 16#0B#),
      2932 => to_slv(opcode_type, 16#0E#),
      2933 => to_slv(opcode_type, 16#08#),
      2934 => to_slv(opcode_type, 16#11#),
      2935 => to_slv(opcode_type, 16#11#),
      2936 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#06#),
      2945 => to_slv(opcode_type, 16#05#),
      2946 => to_slv(opcode_type, 16#06#),
      2947 => to_slv(opcode_type, 16#06#),
      2948 => to_slv(opcode_type, 16#4A#),
      2949 => to_slv(opcode_type, 16#10#),
      2950 => to_slv(opcode_type, 16#06#),
      2951 => to_slv(opcode_type, 16#0E#),
      2952 => to_slv(opcode_type, 16#0F#),
      2953 => to_slv(opcode_type, 16#07#),
      2954 => to_slv(opcode_type, 16#07#),
      2955 => to_slv(opcode_type, 16#08#),
      2956 => to_slv(opcode_type, 16#0C#),
      2957 => to_slv(opcode_type, 16#0B#),
      2958 => to_slv(opcode_type, 16#06#),
      2959 => to_slv(opcode_type, 16#0A#),
      2960 => to_slv(opcode_type, 16#0C#),
      2961 => to_slv(opcode_type, 16#06#),
      2962 => to_slv(opcode_type, 16#07#),
      2963 => to_slv(opcode_type, 16#10#),
      2964 => to_slv(opcode_type, 16#0A#),
      2965 => to_slv(opcode_type, 16#09#),
      2966 => to_slv(opcode_type, 16#0B#),
      2967 => to_slv(opcode_type, 16#0F#),
      2968 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#09#),
      2977 => to_slv(opcode_type, 16#08#),
      2978 => to_slv(opcode_type, 16#07#),
      2979 => to_slv(opcode_type, 16#06#),
      2980 => to_slv(opcode_type, 16#0B#),
      2981 => to_slv(opcode_type, 16#0A#),
      2982 => to_slv(opcode_type, 16#03#),
      2983 => to_slv(opcode_type, 16#C2#),
      2984 => to_slv(opcode_type, 16#05#),
      2985 => to_slv(opcode_type, 16#08#),
      2986 => to_slv(opcode_type, 16#0A#),
      2987 => to_slv(opcode_type, 16#0C#),
      2988 => to_slv(opcode_type, 16#09#),
      2989 => to_slv(opcode_type, 16#03#),
      2990 => to_slv(opcode_type, 16#09#),
      2991 => to_slv(opcode_type, 16#0E#),
      2992 => to_slv(opcode_type, 16#0D#),
      2993 => to_slv(opcode_type, 16#08#),
      2994 => to_slv(opcode_type, 16#09#),
      2995 => to_slv(opcode_type, 16#11#),
      2996 => to_slv(opcode_type, 16#11#),
      2997 => to_slv(opcode_type, 16#07#),
      2998 => to_slv(opcode_type, 16#0A#),
      2999 => to_slv(opcode_type, 16#0B#),
      3000 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#07#),
      3009 => to_slv(opcode_type, 16#03#),
      3010 => to_slv(opcode_type, 16#08#),
      3011 => to_slv(opcode_type, 16#09#),
      3012 => to_slv(opcode_type, 16#0E#),
      3013 => to_slv(opcode_type, 16#0A#),
      3014 => to_slv(opcode_type, 16#09#),
      3015 => to_slv(opcode_type, 16#0B#),
      3016 => to_slv(opcode_type, 16#11#),
      3017 => to_slv(opcode_type, 16#09#),
      3018 => to_slv(opcode_type, 16#06#),
      3019 => to_slv(opcode_type, 16#09#),
      3020 => to_slv(opcode_type, 16#0A#),
      3021 => to_slv(opcode_type, 16#11#),
      3022 => to_slv(opcode_type, 16#08#),
      3023 => to_slv(opcode_type, 16#20#),
      3024 => to_slv(opcode_type, 16#10#),
      3025 => to_slv(opcode_type, 16#09#),
      3026 => to_slv(opcode_type, 16#06#),
      3027 => to_slv(opcode_type, 16#0F#),
      3028 => to_slv(opcode_type, 16#10#),
      3029 => to_slv(opcode_type, 16#08#),
      3030 => to_slv(opcode_type, 16#10#),
      3031 => to_slv(opcode_type, 16#11#),
      3032 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#06#),
      3041 => to_slv(opcode_type, 16#06#),
      3042 => to_slv(opcode_type, 16#09#),
      3043 => to_slv(opcode_type, 16#09#),
      3044 => to_slv(opcode_type, 16#0E#),
      3045 => to_slv(opcode_type, 16#CE#),
      3046 => to_slv(opcode_type, 16#02#),
      3047 => to_slv(opcode_type, 16#0A#),
      3048 => to_slv(opcode_type, 16#03#),
      3049 => to_slv(opcode_type, 16#08#),
      3050 => to_slv(opcode_type, 16#10#),
      3051 => to_slv(opcode_type, 16#0A#),
      3052 => to_slv(opcode_type, 16#06#),
      3053 => to_slv(opcode_type, 16#02#),
      3054 => to_slv(opcode_type, 16#09#),
      3055 => to_slv(opcode_type, 16#11#),
      3056 => to_slv(opcode_type, 16#0F#),
      3057 => to_slv(opcode_type, 16#07#),
      3058 => to_slv(opcode_type, 16#06#),
      3059 => to_slv(opcode_type, 16#0F#),
      3060 => to_slv(opcode_type, 16#11#),
      3061 => to_slv(opcode_type, 16#07#),
      3062 => to_slv(opcode_type, 16#FA#),
      3063 => to_slv(opcode_type, 16#0A#),
      3064 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#08#),
      3073 => to_slv(opcode_type, 16#08#),
      3074 => to_slv(opcode_type, 16#07#),
      3075 => to_slv(opcode_type, 16#08#),
      3076 => to_slv(opcode_type, 16#10#),
      3077 => to_slv(opcode_type, 16#0E#),
      3078 => to_slv(opcode_type, 16#01#),
      3079 => to_slv(opcode_type, 16#0B#),
      3080 => to_slv(opcode_type, 16#05#),
      3081 => to_slv(opcode_type, 16#07#),
      3082 => to_slv(opcode_type, 16#57#),
      3083 => to_slv(opcode_type, 16#10#),
      3084 => to_slv(opcode_type, 16#06#),
      3085 => to_slv(opcode_type, 16#02#),
      3086 => to_slv(opcode_type, 16#09#),
      3087 => to_slv(opcode_type, 16#0D#),
      3088 => to_slv(opcode_type, 16#11#),
      3089 => to_slv(opcode_type, 16#08#),
      3090 => to_slv(opcode_type, 16#06#),
      3091 => to_slv(opcode_type, 16#0F#),
      3092 => to_slv(opcode_type, 16#11#),
      3093 => to_slv(opcode_type, 16#08#),
      3094 => to_slv(opcode_type, 16#0F#),
      3095 => to_slv(opcode_type, 16#B1#),
      3096 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#08#),
      3105 => to_slv(opcode_type, 16#05#),
      3106 => to_slv(opcode_type, 16#09#),
      3107 => to_slv(opcode_type, 16#09#),
      3108 => to_slv(opcode_type, 16#D6#),
      3109 => to_slv(opcode_type, 16#0F#),
      3110 => to_slv(opcode_type, 16#09#),
      3111 => to_slv(opcode_type, 16#0C#),
      3112 => to_slv(opcode_type, 16#0D#),
      3113 => to_slv(opcode_type, 16#08#),
      3114 => to_slv(opcode_type, 16#09#),
      3115 => to_slv(opcode_type, 16#08#),
      3116 => to_slv(opcode_type, 16#11#),
      3117 => to_slv(opcode_type, 16#0A#),
      3118 => to_slv(opcode_type, 16#08#),
      3119 => to_slv(opcode_type, 16#0E#),
      3120 => to_slv(opcode_type, 16#10#),
      3121 => to_slv(opcode_type, 16#06#),
      3122 => to_slv(opcode_type, 16#09#),
      3123 => to_slv(opcode_type, 16#0D#),
      3124 => to_slv(opcode_type, 16#10#),
      3125 => to_slv(opcode_type, 16#07#),
      3126 => to_slv(opcode_type, 16#0C#),
      3127 => to_slv(opcode_type, 16#0E#),
      3128 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#06#),
      3137 => to_slv(opcode_type, 16#06#),
      3138 => to_slv(opcode_type, 16#05#),
      3139 => to_slv(opcode_type, 16#02#),
      3140 => to_slv(opcode_type, 16#BC#),
      3141 => to_slv(opcode_type, 16#02#),
      3142 => to_slv(opcode_type, 16#07#),
      3143 => to_slv(opcode_type, 16#0F#),
      3144 => to_slv(opcode_type, 16#11#),
      3145 => to_slv(opcode_type, 16#07#),
      3146 => to_slv(opcode_type, 16#09#),
      3147 => to_slv(opcode_type, 16#06#),
      3148 => to_slv(opcode_type, 16#5C#),
      3149 => to_slv(opcode_type, 16#10#),
      3150 => to_slv(opcode_type, 16#06#),
      3151 => to_slv(opcode_type, 16#0B#),
      3152 => to_slv(opcode_type, 16#0D#),
      3153 => to_slv(opcode_type, 16#09#),
      3154 => to_slv(opcode_type, 16#07#),
      3155 => to_slv(opcode_type, 16#0E#),
      3156 => to_slv(opcode_type, 16#0F#),
      3157 => to_slv(opcode_type, 16#06#),
      3158 => to_slv(opcode_type, 16#0C#),
      3159 => to_slv(opcode_type, 16#0B#),
      3160 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#06#),
      3169 => to_slv(opcode_type, 16#07#),
      3170 => to_slv(opcode_type, 16#08#),
      3171 => to_slv(opcode_type, 16#07#),
      3172 => to_slv(opcode_type, 16#0F#),
      3173 => to_slv(opcode_type, 16#0E#),
      3174 => to_slv(opcode_type, 16#03#),
      3175 => to_slv(opcode_type, 16#9C#),
      3176 => to_slv(opcode_type, 16#04#),
      3177 => to_slv(opcode_type, 16#05#),
      3178 => to_slv(opcode_type, 16#0E#),
      3179 => to_slv(opcode_type, 16#08#),
      3180 => to_slv(opcode_type, 16#09#),
      3181 => to_slv(opcode_type, 16#02#),
      3182 => to_slv(opcode_type, 16#0F#),
      3183 => to_slv(opcode_type, 16#03#),
      3184 => to_slv(opcode_type, 16#0D#),
      3185 => to_slv(opcode_type, 16#09#),
      3186 => to_slv(opcode_type, 16#07#),
      3187 => to_slv(opcode_type, 16#0C#),
      3188 => to_slv(opcode_type, 16#0C#),
      3189 => to_slv(opcode_type, 16#08#),
      3190 => to_slv(opcode_type, 16#25#),
      3191 => to_slv(opcode_type, 16#0D#),
      3192 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#07#),
      3201 => to_slv(opcode_type, 16#04#),
      3202 => to_slv(opcode_type, 16#06#),
      3203 => to_slv(opcode_type, 16#06#),
      3204 => to_slv(opcode_type, 16#0A#),
      3205 => to_slv(opcode_type, 16#0E#),
      3206 => to_slv(opcode_type, 16#06#),
      3207 => to_slv(opcode_type, 16#3D#),
      3208 => to_slv(opcode_type, 16#0D#),
      3209 => to_slv(opcode_type, 16#09#),
      3210 => to_slv(opcode_type, 16#07#),
      3211 => to_slv(opcode_type, 16#09#),
      3212 => to_slv(opcode_type, 16#AC#),
      3213 => to_slv(opcode_type, 16#0E#),
      3214 => to_slv(opcode_type, 16#08#),
      3215 => to_slv(opcode_type, 16#0E#),
      3216 => to_slv(opcode_type, 16#0F#),
      3217 => to_slv(opcode_type, 16#09#),
      3218 => to_slv(opcode_type, 16#07#),
      3219 => to_slv(opcode_type, 16#0B#),
      3220 => to_slv(opcode_type, 16#0D#),
      3221 => to_slv(opcode_type, 16#08#),
      3222 => to_slv(opcode_type, 16#10#),
      3223 => to_slv(opcode_type, 16#0A#),
      3224 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#07#),
      3233 => to_slv(opcode_type, 16#04#),
      3234 => to_slv(opcode_type, 16#06#),
      3235 => to_slv(opcode_type, 16#06#),
      3236 => to_slv(opcode_type, 16#A0#),
      3237 => to_slv(opcode_type, 16#0D#),
      3238 => to_slv(opcode_type, 16#06#),
      3239 => to_slv(opcode_type, 16#40#),
      3240 => to_slv(opcode_type, 16#0F#),
      3241 => to_slv(opcode_type, 16#06#),
      3242 => to_slv(opcode_type, 16#09#),
      3243 => to_slv(opcode_type, 16#09#),
      3244 => to_slv(opcode_type, 16#0D#),
      3245 => to_slv(opcode_type, 16#0F#),
      3246 => to_slv(opcode_type, 16#07#),
      3247 => to_slv(opcode_type, 16#14#),
      3248 => to_slv(opcode_type, 16#0C#),
      3249 => to_slv(opcode_type, 16#09#),
      3250 => to_slv(opcode_type, 16#06#),
      3251 => to_slv(opcode_type, 16#0A#),
      3252 => to_slv(opcode_type, 16#0E#),
      3253 => to_slv(opcode_type, 16#08#),
      3254 => to_slv(opcode_type, 16#0C#),
      3255 => to_slv(opcode_type, 16#0B#),
      3256 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#06#),
      3265 => to_slv(opcode_type, 16#09#),
      3266 => to_slv(opcode_type, 16#09#),
      3267 => to_slv(opcode_type, 16#01#),
      3268 => to_slv(opcode_type, 16#11#),
      3269 => to_slv(opcode_type, 16#01#),
      3270 => to_slv(opcode_type, 16#0E#),
      3271 => to_slv(opcode_type, 16#08#),
      3272 => to_slv(opcode_type, 16#08#),
      3273 => to_slv(opcode_type, 16#0E#),
      3274 => to_slv(opcode_type, 16#0A#),
      3275 => to_slv(opcode_type, 16#06#),
      3276 => to_slv(opcode_type, 16#10#),
      3277 => to_slv(opcode_type, 16#0F#),
      3278 => to_slv(opcode_type, 16#06#),
      3279 => to_slv(opcode_type, 16#05#),
      3280 => to_slv(opcode_type, 16#01#),
      3281 => to_slv(opcode_type, 16#10#),
      3282 => to_slv(opcode_type, 16#07#),
      3283 => to_slv(opcode_type, 16#01#),
      3284 => to_slv(opcode_type, 16#0E#),
      3285 => to_slv(opcode_type, 16#08#),
      3286 => to_slv(opcode_type, 16#0E#),
      3287 => to_slv(opcode_type, 16#0C#),
      3288 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#07#),
      3297 => to_slv(opcode_type, 16#04#),
      3298 => to_slv(opcode_type, 16#08#),
      3299 => to_slv(opcode_type, 16#08#),
      3300 => to_slv(opcode_type, 16#0B#),
      3301 => to_slv(opcode_type, 16#0D#),
      3302 => to_slv(opcode_type, 16#08#),
      3303 => to_slv(opcode_type, 16#0D#),
      3304 => to_slv(opcode_type, 16#11#),
      3305 => to_slv(opcode_type, 16#08#),
      3306 => to_slv(opcode_type, 16#08#),
      3307 => to_slv(opcode_type, 16#09#),
      3308 => to_slv(opcode_type, 16#0B#),
      3309 => to_slv(opcode_type, 16#11#),
      3310 => to_slv(opcode_type, 16#07#),
      3311 => to_slv(opcode_type, 16#11#),
      3312 => to_slv(opcode_type, 16#0F#),
      3313 => to_slv(opcode_type, 16#09#),
      3314 => to_slv(opcode_type, 16#08#),
      3315 => to_slv(opcode_type, 16#11#),
      3316 => to_slv(opcode_type, 16#10#),
      3317 => to_slv(opcode_type, 16#07#),
      3318 => to_slv(opcode_type, 16#11#),
      3319 => to_slv(opcode_type, 16#11#),
      3320 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#08#),
      3329 => to_slv(opcode_type, 16#04#),
      3330 => to_slv(opcode_type, 16#06#),
      3331 => to_slv(opcode_type, 16#08#),
      3332 => to_slv(opcode_type, 16#0D#),
      3333 => to_slv(opcode_type, 16#0E#),
      3334 => to_slv(opcode_type, 16#08#),
      3335 => to_slv(opcode_type, 16#11#),
      3336 => to_slv(opcode_type, 16#0F#),
      3337 => to_slv(opcode_type, 16#08#),
      3338 => to_slv(opcode_type, 16#08#),
      3339 => to_slv(opcode_type, 16#09#),
      3340 => to_slv(opcode_type, 16#11#),
      3341 => to_slv(opcode_type, 16#CF#),
      3342 => to_slv(opcode_type, 16#09#),
      3343 => to_slv(opcode_type, 16#11#),
      3344 => to_slv(opcode_type, 16#A5#),
      3345 => to_slv(opcode_type, 16#08#),
      3346 => to_slv(opcode_type, 16#09#),
      3347 => to_slv(opcode_type, 16#0E#),
      3348 => to_slv(opcode_type, 16#11#),
      3349 => to_slv(opcode_type, 16#08#),
      3350 => to_slv(opcode_type, 16#0C#),
      3351 => to_slv(opcode_type, 16#11#),
      3352 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#06#),
      3361 => to_slv(opcode_type, 16#09#),
      3362 => to_slv(opcode_type, 16#08#),
      3363 => to_slv(opcode_type, 16#08#),
      3364 => to_slv(opcode_type, 16#11#),
      3365 => to_slv(opcode_type, 16#11#),
      3366 => to_slv(opcode_type, 16#04#),
      3367 => to_slv(opcode_type, 16#76#),
      3368 => to_slv(opcode_type, 16#06#),
      3369 => to_slv(opcode_type, 16#04#),
      3370 => to_slv(opcode_type, 16#0C#),
      3371 => to_slv(opcode_type, 16#05#),
      3372 => to_slv(opcode_type, 16#0F#),
      3373 => to_slv(opcode_type, 16#06#),
      3374 => to_slv(opcode_type, 16#01#),
      3375 => to_slv(opcode_type, 16#09#),
      3376 => to_slv(opcode_type, 16#0C#),
      3377 => to_slv(opcode_type, 16#0E#),
      3378 => to_slv(opcode_type, 16#07#),
      3379 => to_slv(opcode_type, 16#09#),
      3380 => to_slv(opcode_type, 16#11#),
      3381 => to_slv(opcode_type, 16#0F#),
      3382 => to_slv(opcode_type, 16#03#),
      3383 => to_slv(opcode_type, 16#10#),
      3384 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#07#),
      3393 => to_slv(opcode_type, 16#03#),
      3394 => to_slv(opcode_type, 16#06#),
      3395 => to_slv(opcode_type, 16#08#),
      3396 => to_slv(opcode_type, 16#A1#),
      3397 => to_slv(opcode_type, 16#0D#),
      3398 => to_slv(opcode_type, 16#06#),
      3399 => to_slv(opcode_type, 16#0A#),
      3400 => to_slv(opcode_type, 16#0C#),
      3401 => to_slv(opcode_type, 16#06#),
      3402 => to_slv(opcode_type, 16#08#),
      3403 => to_slv(opcode_type, 16#09#),
      3404 => to_slv(opcode_type, 16#6F#),
      3405 => to_slv(opcode_type, 16#0D#),
      3406 => to_slv(opcode_type, 16#09#),
      3407 => to_slv(opcode_type, 16#11#),
      3408 => to_slv(opcode_type, 16#0C#),
      3409 => to_slv(opcode_type, 16#07#),
      3410 => to_slv(opcode_type, 16#09#),
      3411 => to_slv(opcode_type, 16#0E#),
      3412 => to_slv(opcode_type, 16#0A#),
      3413 => to_slv(opcode_type, 16#06#),
      3414 => to_slv(opcode_type, 16#11#),
      3415 => to_slv(opcode_type, 16#5B#),
      3416 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#03#),
      3426 => to_slv(opcode_type, 16#09#),
      3427 => to_slv(opcode_type, 16#06#),
      3428 => to_slv(opcode_type, 16#0F#),
      3429 => to_slv(opcode_type, 16#0A#),
      3430 => to_slv(opcode_type, 16#07#),
      3431 => to_slv(opcode_type, 16#0A#),
      3432 => to_slv(opcode_type, 16#0B#),
      3433 => to_slv(opcode_type, 16#06#),
      3434 => to_slv(opcode_type, 16#06#),
      3435 => to_slv(opcode_type, 16#07#),
      3436 => to_slv(opcode_type, 16#10#),
      3437 => to_slv(opcode_type, 16#51#),
      3438 => to_slv(opcode_type, 16#07#),
      3439 => to_slv(opcode_type, 16#0F#),
      3440 => to_slv(opcode_type, 16#0D#),
      3441 => to_slv(opcode_type, 16#09#),
      3442 => to_slv(opcode_type, 16#08#),
      3443 => to_slv(opcode_type, 16#DF#),
      3444 => to_slv(opcode_type, 16#10#),
      3445 => to_slv(opcode_type, 16#08#),
      3446 => to_slv(opcode_type, 16#0A#),
      3447 => to_slv(opcode_type, 16#0B#),
      3448 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#08#),
      3457 => to_slv(opcode_type, 16#06#),
      3458 => to_slv(opcode_type, 16#02#),
      3459 => to_slv(opcode_type, 16#08#),
      3460 => to_slv(opcode_type, 16#0B#),
      3461 => to_slv(opcode_type, 16#40#),
      3462 => to_slv(opcode_type, 16#09#),
      3463 => to_slv(opcode_type, 16#09#),
      3464 => to_slv(opcode_type, 16#DE#),
      3465 => to_slv(opcode_type, 16#0F#),
      3466 => to_slv(opcode_type, 16#08#),
      3467 => to_slv(opcode_type, 16#0B#),
      3468 => to_slv(opcode_type, 16#11#),
      3469 => to_slv(opcode_type, 16#09#),
      3470 => to_slv(opcode_type, 16#03#),
      3471 => to_slv(opcode_type, 16#04#),
      3472 => to_slv(opcode_type, 16#0B#),
      3473 => to_slv(opcode_type, 16#07#),
      3474 => to_slv(opcode_type, 16#06#),
      3475 => to_slv(opcode_type, 16#0A#),
      3476 => to_slv(opcode_type, 16#0D#),
      3477 => to_slv(opcode_type, 16#09#),
      3478 => to_slv(opcode_type, 16#10#),
      3479 => to_slv(opcode_type, 16#0D#),
      3480 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#09#),
      3489 => to_slv(opcode_type, 16#03#),
      3490 => to_slv(opcode_type, 16#06#),
      3491 => to_slv(opcode_type, 16#06#),
      3492 => to_slv(opcode_type, 16#4B#),
      3493 => to_slv(opcode_type, 16#0D#),
      3494 => to_slv(opcode_type, 16#09#),
      3495 => to_slv(opcode_type, 16#11#),
      3496 => to_slv(opcode_type, 16#0C#),
      3497 => to_slv(opcode_type, 16#07#),
      3498 => to_slv(opcode_type, 16#08#),
      3499 => to_slv(opcode_type, 16#09#),
      3500 => to_slv(opcode_type, 16#0C#),
      3501 => to_slv(opcode_type, 16#0D#),
      3502 => to_slv(opcode_type, 16#06#),
      3503 => to_slv(opcode_type, 16#0C#),
      3504 => to_slv(opcode_type, 16#0E#),
      3505 => to_slv(opcode_type, 16#09#),
      3506 => to_slv(opcode_type, 16#09#),
      3507 => to_slv(opcode_type, 16#0A#),
      3508 => to_slv(opcode_type, 16#0D#),
      3509 => to_slv(opcode_type, 16#09#),
      3510 => to_slv(opcode_type, 16#0E#),
      3511 => to_slv(opcode_type, 16#0A#),
      3512 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#09#),
      3521 => to_slv(opcode_type, 16#04#),
      3522 => to_slv(opcode_type, 16#09#),
      3523 => to_slv(opcode_type, 16#09#),
      3524 => to_slv(opcode_type, 16#11#),
      3525 => to_slv(opcode_type, 16#11#),
      3526 => to_slv(opcode_type, 16#08#),
      3527 => to_slv(opcode_type, 16#3C#),
      3528 => to_slv(opcode_type, 16#0E#),
      3529 => to_slv(opcode_type, 16#07#),
      3530 => to_slv(opcode_type, 16#09#),
      3531 => to_slv(opcode_type, 16#06#),
      3532 => to_slv(opcode_type, 16#0C#),
      3533 => to_slv(opcode_type, 16#0F#),
      3534 => to_slv(opcode_type, 16#08#),
      3535 => to_slv(opcode_type, 16#0C#),
      3536 => to_slv(opcode_type, 16#0E#),
      3537 => to_slv(opcode_type, 16#07#),
      3538 => to_slv(opcode_type, 16#09#),
      3539 => to_slv(opcode_type, 16#0C#),
      3540 => to_slv(opcode_type, 16#0F#),
      3541 => to_slv(opcode_type, 16#07#),
      3542 => to_slv(opcode_type, 16#0C#),
      3543 => to_slv(opcode_type, 16#10#),
      3544 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#08#),
      3553 => to_slv(opcode_type, 16#09#),
      3554 => to_slv(opcode_type, 16#05#),
      3555 => to_slv(opcode_type, 16#05#),
      3556 => to_slv(opcode_type, 16#0A#),
      3557 => to_slv(opcode_type, 16#04#),
      3558 => to_slv(opcode_type, 16#09#),
      3559 => to_slv(opcode_type, 16#0E#),
      3560 => to_slv(opcode_type, 16#0D#),
      3561 => to_slv(opcode_type, 16#06#),
      3562 => to_slv(opcode_type, 16#08#),
      3563 => to_slv(opcode_type, 16#06#),
      3564 => to_slv(opcode_type, 16#11#),
      3565 => to_slv(opcode_type, 16#11#),
      3566 => to_slv(opcode_type, 16#06#),
      3567 => to_slv(opcode_type, 16#0E#),
      3568 => to_slv(opcode_type, 16#0D#),
      3569 => to_slv(opcode_type, 16#09#),
      3570 => to_slv(opcode_type, 16#07#),
      3571 => to_slv(opcode_type, 16#10#),
      3572 => to_slv(opcode_type, 16#0B#),
      3573 => to_slv(opcode_type, 16#07#),
      3574 => to_slv(opcode_type, 16#11#),
      3575 => to_slv(opcode_type, 16#0D#),
      3576 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#06#),
      3585 => to_slv(opcode_type, 16#02#),
      3586 => to_slv(opcode_type, 16#07#),
      3587 => to_slv(opcode_type, 16#07#),
      3588 => to_slv(opcode_type, 16#0C#),
      3589 => to_slv(opcode_type, 16#0B#),
      3590 => to_slv(opcode_type, 16#08#),
      3591 => to_slv(opcode_type, 16#10#),
      3592 => to_slv(opcode_type, 16#0F#),
      3593 => to_slv(opcode_type, 16#06#),
      3594 => to_slv(opcode_type, 16#07#),
      3595 => to_slv(opcode_type, 16#06#),
      3596 => to_slv(opcode_type, 16#10#),
      3597 => to_slv(opcode_type, 16#0F#),
      3598 => to_slv(opcode_type, 16#09#),
      3599 => to_slv(opcode_type, 16#0A#),
      3600 => to_slv(opcode_type, 16#0A#),
      3601 => to_slv(opcode_type, 16#08#),
      3602 => to_slv(opcode_type, 16#09#),
      3603 => to_slv(opcode_type, 16#F5#),
      3604 => to_slv(opcode_type, 16#0D#),
      3605 => to_slv(opcode_type, 16#06#),
      3606 => to_slv(opcode_type, 16#FA#),
      3607 => to_slv(opcode_type, 16#0B#),
      3608 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#07#),
      3617 => to_slv(opcode_type, 16#01#),
      3618 => to_slv(opcode_type, 16#09#),
      3619 => to_slv(opcode_type, 16#08#),
      3620 => to_slv(opcode_type, 16#90#),
      3621 => to_slv(opcode_type, 16#11#),
      3622 => to_slv(opcode_type, 16#07#),
      3623 => to_slv(opcode_type, 16#0A#),
      3624 => to_slv(opcode_type, 16#10#),
      3625 => to_slv(opcode_type, 16#09#),
      3626 => to_slv(opcode_type, 16#07#),
      3627 => to_slv(opcode_type, 16#08#),
      3628 => to_slv(opcode_type, 16#4B#),
      3629 => to_slv(opcode_type, 16#11#),
      3630 => to_slv(opcode_type, 16#06#),
      3631 => to_slv(opcode_type, 16#0E#),
      3632 => to_slv(opcode_type, 16#2B#),
      3633 => to_slv(opcode_type, 16#07#),
      3634 => to_slv(opcode_type, 16#06#),
      3635 => to_slv(opcode_type, 16#0F#),
      3636 => to_slv(opcode_type, 16#F4#),
      3637 => to_slv(opcode_type, 16#09#),
      3638 => to_slv(opcode_type, 16#11#),
      3639 => to_slv(opcode_type, 16#0E#),
      3640 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#06#),
      3649 => to_slv(opcode_type, 16#06#),
      3650 => to_slv(opcode_type, 16#04#),
      3651 => to_slv(opcode_type, 16#04#),
      3652 => to_slv(opcode_type, 16#B5#),
      3653 => to_slv(opcode_type, 16#05#),
      3654 => to_slv(opcode_type, 16#07#),
      3655 => to_slv(opcode_type, 16#0F#),
      3656 => to_slv(opcode_type, 16#0E#),
      3657 => to_slv(opcode_type, 16#09#),
      3658 => to_slv(opcode_type, 16#06#),
      3659 => to_slv(opcode_type, 16#09#),
      3660 => to_slv(opcode_type, 16#10#),
      3661 => to_slv(opcode_type, 16#11#),
      3662 => to_slv(opcode_type, 16#07#),
      3663 => to_slv(opcode_type, 16#AD#),
      3664 => to_slv(opcode_type, 16#0B#),
      3665 => to_slv(opcode_type, 16#08#),
      3666 => to_slv(opcode_type, 16#09#),
      3667 => to_slv(opcode_type, 16#0D#),
      3668 => to_slv(opcode_type, 16#B6#),
      3669 => to_slv(opcode_type, 16#07#),
      3670 => to_slv(opcode_type, 16#DD#),
      3671 => to_slv(opcode_type, 16#0A#),
      3672 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#09#),
      3681 => to_slv(opcode_type, 16#08#),
      3682 => to_slv(opcode_type, 16#05#),
      3683 => to_slv(opcode_type, 16#01#),
      3684 => to_slv(opcode_type, 16#0E#),
      3685 => to_slv(opcode_type, 16#08#),
      3686 => to_slv(opcode_type, 16#07#),
      3687 => to_slv(opcode_type, 16#0E#),
      3688 => to_slv(opcode_type, 16#0A#),
      3689 => to_slv(opcode_type, 16#02#),
      3690 => to_slv(opcode_type, 16#0E#),
      3691 => to_slv(opcode_type, 16#06#),
      3692 => to_slv(opcode_type, 16#07#),
      3693 => to_slv(opcode_type, 16#06#),
      3694 => to_slv(opcode_type, 16#11#),
      3695 => to_slv(opcode_type, 16#D6#),
      3696 => to_slv(opcode_type, 16#08#),
      3697 => to_slv(opcode_type, 16#0B#),
      3698 => to_slv(opcode_type, 16#10#),
      3699 => to_slv(opcode_type, 16#08#),
      3700 => to_slv(opcode_type, 16#03#),
      3701 => to_slv(opcode_type, 16#0F#),
      3702 => to_slv(opcode_type, 16#02#),
      3703 => to_slv(opcode_type, 16#0B#),
      3704 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#09#),
      3713 => to_slv(opcode_type, 16#09#),
      3714 => to_slv(opcode_type, 16#04#),
      3715 => to_slv(opcode_type, 16#03#),
      3716 => to_slv(opcode_type, 16#0F#),
      3717 => to_slv(opcode_type, 16#05#),
      3718 => to_slv(opcode_type, 16#09#),
      3719 => to_slv(opcode_type, 16#0D#),
      3720 => to_slv(opcode_type, 16#0A#),
      3721 => to_slv(opcode_type, 16#08#),
      3722 => to_slv(opcode_type, 16#08#),
      3723 => to_slv(opcode_type, 16#07#),
      3724 => to_slv(opcode_type, 16#0E#),
      3725 => to_slv(opcode_type, 16#11#),
      3726 => to_slv(opcode_type, 16#08#),
      3727 => to_slv(opcode_type, 16#10#),
      3728 => to_slv(opcode_type, 16#11#),
      3729 => to_slv(opcode_type, 16#06#),
      3730 => to_slv(opcode_type, 16#09#),
      3731 => to_slv(opcode_type, 16#0A#),
      3732 => to_slv(opcode_type, 16#44#),
      3733 => to_slv(opcode_type, 16#07#),
      3734 => to_slv(opcode_type, 16#11#),
      3735 => to_slv(opcode_type, 16#0B#),
      3736 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#08#),
      3745 => to_slv(opcode_type, 16#06#),
      3746 => to_slv(opcode_type, 16#02#),
      3747 => to_slv(opcode_type, 16#07#),
      3748 => to_slv(opcode_type, 16#0E#),
      3749 => to_slv(opcode_type, 16#0A#),
      3750 => to_slv(opcode_type, 16#08#),
      3751 => to_slv(opcode_type, 16#08#),
      3752 => to_slv(opcode_type, 16#0D#),
      3753 => to_slv(opcode_type, 16#6E#),
      3754 => to_slv(opcode_type, 16#01#),
      3755 => to_slv(opcode_type, 16#0A#),
      3756 => to_slv(opcode_type, 16#08#),
      3757 => to_slv(opcode_type, 16#06#),
      3758 => to_slv(opcode_type, 16#08#),
      3759 => to_slv(opcode_type, 16#10#),
      3760 => to_slv(opcode_type, 16#11#),
      3761 => to_slv(opcode_type, 16#09#),
      3762 => to_slv(opcode_type, 16#11#),
      3763 => to_slv(opcode_type, 16#0A#),
      3764 => to_slv(opcode_type, 16#05#),
      3765 => to_slv(opcode_type, 16#09#),
      3766 => to_slv(opcode_type, 16#0A#),
      3767 => to_slv(opcode_type, 16#0C#),
      3768 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#07#),
      3777 => to_slv(opcode_type, 16#01#),
      3778 => to_slv(opcode_type, 16#09#),
      3779 => to_slv(opcode_type, 16#06#),
      3780 => to_slv(opcode_type, 16#11#),
      3781 => to_slv(opcode_type, 16#0E#),
      3782 => to_slv(opcode_type, 16#08#),
      3783 => to_slv(opcode_type, 16#0D#),
      3784 => to_slv(opcode_type, 16#0A#),
      3785 => to_slv(opcode_type, 16#07#),
      3786 => to_slv(opcode_type, 16#08#),
      3787 => to_slv(opcode_type, 16#06#),
      3788 => to_slv(opcode_type, 16#0D#),
      3789 => to_slv(opcode_type, 16#0F#),
      3790 => to_slv(opcode_type, 16#07#),
      3791 => to_slv(opcode_type, 16#0F#),
      3792 => to_slv(opcode_type, 16#0B#),
      3793 => to_slv(opcode_type, 16#07#),
      3794 => to_slv(opcode_type, 16#08#),
      3795 => to_slv(opcode_type, 16#0B#),
      3796 => to_slv(opcode_type, 16#0A#),
      3797 => to_slv(opcode_type, 16#09#),
      3798 => to_slv(opcode_type, 16#10#),
      3799 => to_slv(opcode_type, 16#0D#),
      3800 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#08#),
      3809 => to_slv(opcode_type, 16#02#),
      3810 => to_slv(opcode_type, 16#09#),
      3811 => to_slv(opcode_type, 16#08#),
      3812 => to_slv(opcode_type, 16#11#),
      3813 => to_slv(opcode_type, 16#0F#),
      3814 => to_slv(opcode_type, 16#07#),
      3815 => to_slv(opcode_type, 16#10#),
      3816 => to_slv(opcode_type, 16#0A#),
      3817 => to_slv(opcode_type, 16#09#),
      3818 => to_slv(opcode_type, 16#08#),
      3819 => to_slv(opcode_type, 16#06#),
      3820 => to_slv(opcode_type, 16#0B#),
      3821 => to_slv(opcode_type, 16#0E#),
      3822 => to_slv(opcode_type, 16#06#),
      3823 => to_slv(opcode_type, 16#0A#),
      3824 => to_slv(opcode_type, 16#0A#),
      3825 => to_slv(opcode_type, 16#07#),
      3826 => to_slv(opcode_type, 16#06#),
      3827 => to_slv(opcode_type, 16#0D#),
      3828 => to_slv(opcode_type, 16#4E#),
      3829 => to_slv(opcode_type, 16#09#),
      3830 => to_slv(opcode_type, 16#10#),
      3831 => to_slv(opcode_type, 16#68#),
      3832 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#07#),
      3841 => to_slv(opcode_type, 16#04#),
      3842 => to_slv(opcode_type, 16#06#),
      3843 => to_slv(opcode_type, 16#09#),
      3844 => to_slv(opcode_type, 16#28#),
      3845 => to_slv(opcode_type, 16#11#),
      3846 => to_slv(opcode_type, 16#07#),
      3847 => to_slv(opcode_type, 16#0B#),
      3848 => to_slv(opcode_type, 16#17#),
      3849 => to_slv(opcode_type, 16#08#),
      3850 => to_slv(opcode_type, 16#09#),
      3851 => to_slv(opcode_type, 16#07#),
      3852 => to_slv(opcode_type, 16#0E#),
      3853 => to_slv(opcode_type, 16#10#),
      3854 => to_slv(opcode_type, 16#07#),
      3855 => to_slv(opcode_type, 16#0B#),
      3856 => to_slv(opcode_type, 16#0E#),
      3857 => to_slv(opcode_type, 16#07#),
      3858 => to_slv(opcode_type, 16#06#),
      3859 => to_slv(opcode_type, 16#0E#),
      3860 => to_slv(opcode_type, 16#24#),
      3861 => to_slv(opcode_type, 16#08#),
      3862 => to_slv(opcode_type, 16#10#),
      3863 => to_slv(opcode_type, 16#0B#),
      3864 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#09#),
      3873 => to_slv(opcode_type, 16#09#),
      3874 => to_slv(opcode_type, 16#09#),
      3875 => to_slv(opcode_type, 16#04#),
      3876 => to_slv(opcode_type, 16#57#),
      3877 => to_slv(opcode_type, 16#02#),
      3878 => to_slv(opcode_type, 16#0A#),
      3879 => to_slv(opcode_type, 16#09#),
      3880 => to_slv(opcode_type, 16#07#),
      3881 => to_slv(opcode_type, 16#10#),
      3882 => to_slv(opcode_type, 16#11#),
      3883 => to_slv(opcode_type, 16#06#),
      3884 => to_slv(opcode_type, 16#0F#),
      3885 => to_slv(opcode_type, 16#0B#),
      3886 => to_slv(opcode_type, 16#07#),
      3887 => to_slv(opcode_type, 16#03#),
      3888 => to_slv(opcode_type, 16#08#),
      3889 => to_slv(opcode_type, 16#11#),
      3890 => to_slv(opcode_type, 16#0F#),
      3891 => to_slv(opcode_type, 16#09#),
      3892 => to_slv(opcode_type, 16#09#),
      3893 => to_slv(opcode_type, 16#11#),
      3894 => to_slv(opcode_type, 16#0A#),
      3895 => to_slv(opcode_type, 16#0F#),
      3896 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#08#),
      3905 => to_slv(opcode_type, 16#09#),
      3906 => to_slv(opcode_type, 16#03#),
      3907 => to_slv(opcode_type, 16#03#),
      3908 => to_slv(opcode_type, 16#0B#),
      3909 => to_slv(opcode_type, 16#01#),
      3910 => to_slv(opcode_type, 16#09#),
      3911 => to_slv(opcode_type, 16#0E#),
      3912 => to_slv(opcode_type, 16#0A#),
      3913 => to_slv(opcode_type, 16#08#),
      3914 => to_slv(opcode_type, 16#08#),
      3915 => to_slv(opcode_type, 16#09#),
      3916 => to_slv(opcode_type, 16#11#),
      3917 => to_slv(opcode_type, 16#0E#),
      3918 => to_slv(opcode_type, 16#06#),
      3919 => to_slv(opcode_type, 16#0D#),
      3920 => to_slv(opcode_type, 16#10#),
      3921 => to_slv(opcode_type, 16#06#),
      3922 => to_slv(opcode_type, 16#09#),
      3923 => to_slv(opcode_type, 16#0F#),
      3924 => to_slv(opcode_type, 16#7C#),
      3925 => to_slv(opcode_type, 16#08#),
      3926 => to_slv(opcode_type, 16#0B#),
      3927 => to_slv(opcode_type, 16#0E#),
      3928 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#08#),
      3937 => to_slv(opcode_type, 16#03#),
      3938 => to_slv(opcode_type, 16#08#),
      3939 => to_slv(opcode_type, 16#06#),
      3940 => to_slv(opcode_type, 16#0F#),
      3941 => to_slv(opcode_type, 16#0A#),
      3942 => to_slv(opcode_type, 16#06#),
      3943 => to_slv(opcode_type, 16#0E#),
      3944 => to_slv(opcode_type, 16#6C#),
      3945 => to_slv(opcode_type, 16#08#),
      3946 => to_slv(opcode_type, 16#08#),
      3947 => to_slv(opcode_type, 16#06#),
      3948 => to_slv(opcode_type, 16#0B#),
      3949 => to_slv(opcode_type, 16#0F#),
      3950 => to_slv(opcode_type, 16#08#),
      3951 => to_slv(opcode_type, 16#0B#),
      3952 => to_slv(opcode_type, 16#11#),
      3953 => to_slv(opcode_type, 16#06#),
      3954 => to_slv(opcode_type, 16#08#),
      3955 => to_slv(opcode_type, 16#0F#),
      3956 => to_slv(opcode_type, 16#0B#),
      3957 => to_slv(opcode_type, 16#06#),
      3958 => to_slv(opcode_type, 16#0C#),
      3959 => to_slv(opcode_type, 16#0E#),
      3960 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#08#),
      3969 => to_slv(opcode_type, 16#01#),
      3970 => to_slv(opcode_type, 16#08#),
      3971 => to_slv(opcode_type, 16#07#),
      3972 => to_slv(opcode_type, 16#11#),
      3973 => to_slv(opcode_type, 16#0E#),
      3974 => to_slv(opcode_type, 16#06#),
      3975 => to_slv(opcode_type, 16#0C#),
      3976 => to_slv(opcode_type, 16#AD#),
      3977 => to_slv(opcode_type, 16#07#),
      3978 => to_slv(opcode_type, 16#06#),
      3979 => to_slv(opcode_type, 16#07#),
      3980 => to_slv(opcode_type, 16#10#),
      3981 => to_slv(opcode_type, 16#0D#),
      3982 => to_slv(opcode_type, 16#06#),
      3983 => to_slv(opcode_type, 16#11#),
      3984 => to_slv(opcode_type, 16#0A#),
      3985 => to_slv(opcode_type, 16#08#),
      3986 => to_slv(opcode_type, 16#08#),
      3987 => to_slv(opcode_type, 16#10#),
      3988 => to_slv(opcode_type, 16#0E#),
      3989 => to_slv(opcode_type, 16#09#),
      3990 => to_slv(opcode_type, 16#10#),
      3991 => to_slv(opcode_type, 16#0C#),
      3992 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#06#),
      4001 => to_slv(opcode_type, 16#03#),
      4002 => to_slv(opcode_type, 16#08#),
      4003 => to_slv(opcode_type, 16#09#),
      4004 => to_slv(opcode_type, 16#0B#),
      4005 => to_slv(opcode_type, 16#0C#),
      4006 => to_slv(opcode_type, 16#08#),
      4007 => to_slv(opcode_type, 16#0D#),
      4008 => to_slv(opcode_type, 16#0D#),
      4009 => to_slv(opcode_type, 16#07#),
      4010 => to_slv(opcode_type, 16#09#),
      4011 => to_slv(opcode_type, 16#07#),
      4012 => to_slv(opcode_type, 16#10#),
      4013 => to_slv(opcode_type, 16#0E#),
      4014 => to_slv(opcode_type, 16#07#),
      4015 => to_slv(opcode_type, 16#10#),
      4016 => to_slv(opcode_type, 16#10#),
      4017 => to_slv(opcode_type, 16#08#),
      4018 => to_slv(opcode_type, 16#08#),
      4019 => to_slv(opcode_type, 16#0A#),
      4020 => to_slv(opcode_type, 16#0C#),
      4021 => to_slv(opcode_type, 16#06#),
      4022 => to_slv(opcode_type, 16#11#),
      4023 => to_slv(opcode_type, 16#0D#),
      4024 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#06#),
      4033 => to_slv(opcode_type, 16#03#),
      4034 => to_slv(opcode_type, 16#09#),
      4035 => to_slv(opcode_type, 16#07#),
      4036 => to_slv(opcode_type, 16#0E#),
      4037 => to_slv(opcode_type, 16#0A#),
      4038 => to_slv(opcode_type, 16#08#),
      4039 => to_slv(opcode_type, 16#0A#),
      4040 => to_slv(opcode_type, 16#0D#),
      4041 => to_slv(opcode_type, 16#06#),
      4042 => to_slv(opcode_type, 16#06#),
      4043 => to_slv(opcode_type, 16#07#),
      4044 => to_slv(opcode_type, 16#0E#),
      4045 => to_slv(opcode_type, 16#0A#),
      4046 => to_slv(opcode_type, 16#08#),
      4047 => to_slv(opcode_type, 16#0A#),
      4048 => to_slv(opcode_type, 16#0D#),
      4049 => to_slv(opcode_type, 16#09#),
      4050 => to_slv(opcode_type, 16#06#),
      4051 => to_slv(opcode_type, 16#0E#),
      4052 => to_slv(opcode_type, 16#10#),
      4053 => to_slv(opcode_type, 16#09#),
      4054 => to_slv(opcode_type, 16#0D#),
      4055 => to_slv(opcode_type, 16#0A#),
      4056 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#09#),
      4065 => to_slv(opcode_type, 16#07#),
      4066 => to_slv(opcode_type, 16#08#),
      4067 => to_slv(opcode_type, 16#04#),
      4068 => to_slv(opcode_type, 16#10#),
      4069 => to_slv(opcode_type, 16#08#),
      4070 => to_slv(opcode_type, 16#0D#),
      4071 => to_slv(opcode_type, 16#0A#),
      4072 => to_slv(opcode_type, 16#04#),
      4073 => to_slv(opcode_type, 16#06#),
      4074 => to_slv(opcode_type, 16#11#),
      4075 => to_slv(opcode_type, 16#0A#),
      4076 => to_slv(opcode_type, 16#07#),
      4077 => to_slv(opcode_type, 16#08#),
      4078 => to_slv(opcode_type, 16#06#),
      4079 => to_slv(opcode_type, 16#10#),
      4080 => to_slv(opcode_type, 16#0D#),
      4081 => to_slv(opcode_type, 16#03#),
      4082 => to_slv(opcode_type, 16#EE#),
      4083 => to_slv(opcode_type, 16#06#),
      4084 => to_slv(opcode_type, 16#01#),
      4085 => to_slv(opcode_type, 16#0A#),
      4086 => to_slv(opcode_type, 16#05#),
      4087 => to_slv(opcode_type, 16#CA#),
      4088 to 4095 => (others => '0')
  ),

    -- Bin `25`...
    24 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#06#),
      1 => to_slv(opcode_type, 16#09#),
      2 => to_slv(opcode_type, 16#07#),
      3 => to_slv(opcode_type, 16#07#),
      4 => to_slv(opcode_type, 16#11#),
      5 => to_slv(opcode_type, 16#0D#),
      6 => to_slv(opcode_type, 16#05#),
      7 => to_slv(opcode_type, 16#0C#),
      8 => to_slv(opcode_type, 16#03#),
      9 => to_slv(opcode_type, 16#03#),
      10 => to_slv(opcode_type, 16#10#),
      11 => to_slv(opcode_type, 16#08#),
      12 => to_slv(opcode_type, 16#07#),
      13 => to_slv(opcode_type, 16#03#),
      14 => to_slv(opcode_type, 16#10#),
      15 => to_slv(opcode_type, 16#07#),
      16 => to_slv(opcode_type, 16#0B#),
      17 => to_slv(opcode_type, 16#0D#),
      18 => to_slv(opcode_type, 16#06#),
      19 => to_slv(opcode_type, 16#07#),
      20 => to_slv(opcode_type, 16#10#),
      21 => to_slv(opcode_type, 16#0F#),
      22 => to_slv(opcode_type, 16#07#),
      23 => to_slv(opcode_type, 16#0E#),
      24 => to_slv(opcode_type, 16#0D#),
      25 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#09#),
      33 => to_slv(opcode_type, 16#06#),
      34 => to_slv(opcode_type, 16#05#),
      35 => to_slv(opcode_type, 16#05#),
      36 => to_slv(opcode_type, 16#0D#),
      37 => to_slv(opcode_type, 16#07#),
      38 => to_slv(opcode_type, 16#04#),
      39 => to_slv(opcode_type, 16#0F#),
      40 => to_slv(opcode_type, 16#02#),
      41 => to_slv(opcode_type, 16#0E#),
      42 => to_slv(opcode_type, 16#09#),
      43 => to_slv(opcode_type, 16#08#),
      44 => to_slv(opcode_type, 16#08#),
      45 => to_slv(opcode_type, 16#0B#),
      46 => to_slv(opcode_type, 16#0F#),
      47 => to_slv(opcode_type, 16#08#),
      48 => to_slv(opcode_type, 16#0C#),
      49 => to_slv(opcode_type, 16#0A#),
      50 => to_slv(opcode_type, 16#08#),
      51 => to_slv(opcode_type, 16#06#),
      52 => to_slv(opcode_type, 16#10#),
      53 => to_slv(opcode_type, 16#E2#),
      54 => to_slv(opcode_type, 16#09#),
      55 => to_slv(opcode_type, 16#11#),
      56 => to_slv(opcode_type, 16#0B#),
      57 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#08#),
      65 => to_slv(opcode_type, 16#09#),
      66 => to_slv(opcode_type, 16#05#),
      67 => to_slv(opcode_type, 16#03#),
      68 => to_slv(opcode_type, 16#0D#),
      69 => to_slv(opcode_type, 16#06#),
      70 => to_slv(opcode_type, 16#08#),
      71 => to_slv(opcode_type, 16#0C#),
      72 => to_slv(opcode_type, 16#0A#),
      73 => to_slv(opcode_type, 16#02#),
      74 => to_slv(opcode_type, 16#0D#),
      75 => to_slv(opcode_type, 16#09#),
      76 => to_slv(opcode_type, 16#09#),
      77 => to_slv(opcode_type, 16#08#),
      78 => to_slv(opcode_type, 16#11#),
      79 => to_slv(opcode_type, 16#0A#),
      80 => to_slv(opcode_type, 16#01#),
      81 => to_slv(opcode_type, 16#0A#),
      82 => to_slv(opcode_type, 16#09#),
      83 => to_slv(opcode_type, 16#08#),
      84 => to_slv(opcode_type, 16#0B#),
      85 => to_slv(opcode_type, 16#0F#),
      86 => to_slv(opcode_type, 16#06#),
      87 => to_slv(opcode_type, 16#0F#),
      88 => to_slv(opcode_type, 16#0A#),
      89 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#08#),
      97 => to_slv(opcode_type, 16#09#),
      98 => to_slv(opcode_type, 16#04#),
      99 => to_slv(opcode_type, 16#02#),
      100 => to_slv(opcode_type, 16#0D#),
      101 => to_slv(opcode_type, 16#09#),
      102 => to_slv(opcode_type, 16#04#),
      103 => to_slv(opcode_type, 16#10#),
      104 => to_slv(opcode_type, 16#01#),
      105 => to_slv(opcode_type, 16#0C#),
      106 => to_slv(opcode_type, 16#06#),
      107 => to_slv(opcode_type, 16#09#),
      108 => to_slv(opcode_type, 16#07#),
      109 => to_slv(opcode_type, 16#11#),
      110 => to_slv(opcode_type, 16#0F#),
      111 => to_slv(opcode_type, 16#06#),
      112 => to_slv(opcode_type, 16#0F#),
      113 => to_slv(opcode_type, 16#10#),
      114 => to_slv(opcode_type, 16#06#),
      115 => to_slv(opcode_type, 16#07#),
      116 => to_slv(opcode_type, 16#0D#),
      117 => to_slv(opcode_type, 16#0E#),
      118 => to_slv(opcode_type, 16#08#),
      119 => to_slv(opcode_type, 16#0D#),
      120 => to_slv(opcode_type, 16#0B#),
      121 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#06#),
      129 => to_slv(opcode_type, 16#09#),
      130 => to_slv(opcode_type, 16#04#),
      131 => to_slv(opcode_type, 16#09#),
      132 => to_slv(opcode_type, 16#11#),
      133 => to_slv(opcode_type, 16#11#),
      134 => to_slv(opcode_type, 16#08#),
      135 => to_slv(opcode_type, 16#01#),
      136 => to_slv(opcode_type, 16#0C#),
      137 => to_slv(opcode_type, 16#05#),
      138 => to_slv(opcode_type, 16#0D#),
      139 => to_slv(opcode_type, 16#08#),
      140 => to_slv(opcode_type, 16#08#),
      141 => to_slv(opcode_type, 16#01#),
      142 => to_slv(opcode_type, 16#10#),
      143 => to_slv(opcode_type, 16#09#),
      144 => to_slv(opcode_type, 16#0C#),
      145 => to_slv(opcode_type, 16#11#),
      146 => to_slv(opcode_type, 16#07#),
      147 => to_slv(opcode_type, 16#06#),
      148 => to_slv(opcode_type, 16#10#),
      149 => to_slv(opcode_type, 16#10#),
      150 => to_slv(opcode_type, 16#07#),
      151 => to_slv(opcode_type, 16#0D#),
      152 => to_slv(opcode_type, 16#0D#),
      153 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#08#),
      161 => to_slv(opcode_type, 16#07#),
      162 => to_slv(opcode_type, 16#07#),
      163 => to_slv(opcode_type, 16#06#),
      164 => to_slv(opcode_type, 16#0F#),
      165 => to_slv(opcode_type, 16#0A#),
      166 => to_slv(opcode_type, 16#06#),
      167 => to_slv(opcode_type, 16#10#),
      168 => to_slv(opcode_type, 16#0E#),
      169 => to_slv(opcode_type, 16#03#),
      170 => to_slv(opcode_type, 16#02#),
      171 => to_slv(opcode_type, 16#11#),
      172 => to_slv(opcode_type, 16#07#),
      173 => to_slv(opcode_type, 16#06#),
      174 => to_slv(opcode_type, 16#07#),
      175 => to_slv(opcode_type, 16#10#),
      176 => to_slv(opcode_type, 16#0F#),
      177 => to_slv(opcode_type, 16#06#),
      178 => to_slv(opcode_type, 16#0E#),
      179 => to_slv(opcode_type, 16#0F#),
      180 => to_slv(opcode_type, 16#06#),
      181 => to_slv(opcode_type, 16#02#),
      182 => to_slv(opcode_type, 16#0B#),
      183 => to_slv(opcode_type, 16#02#),
      184 => to_slv(opcode_type, 16#0B#),
      185 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#09#),
      193 => to_slv(opcode_type, 16#08#),
      194 => to_slv(opcode_type, 16#08#),
      195 => to_slv(opcode_type, 16#08#),
      196 => to_slv(opcode_type, 16#0D#),
      197 => to_slv(opcode_type, 16#0F#),
      198 => to_slv(opcode_type, 16#06#),
      199 => to_slv(opcode_type, 16#11#),
      200 => to_slv(opcode_type, 16#0A#),
      201 => to_slv(opcode_type, 16#04#),
      202 => to_slv(opcode_type, 16#07#),
      203 => to_slv(opcode_type, 16#0A#),
      204 => to_slv(opcode_type, 16#0F#),
      205 => to_slv(opcode_type, 16#06#),
      206 => to_slv(opcode_type, 16#01#),
      207 => to_slv(opcode_type, 16#08#),
      208 => to_slv(opcode_type, 16#0F#),
      209 => to_slv(opcode_type, 16#0F#),
      210 => to_slv(opcode_type, 16#07#),
      211 => to_slv(opcode_type, 16#08#),
      212 => to_slv(opcode_type, 16#0D#),
      213 => to_slv(opcode_type, 16#11#),
      214 => to_slv(opcode_type, 16#06#),
      215 => to_slv(opcode_type, 16#0B#),
      216 => to_slv(opcode_type, 16#11#),
      217 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#09#),
      225 => to_slv(opcode_type, 16#09#),
      226 => to_slv(opcode_type, 16#01#),
      227 => to_slv(opcode_type, 16#07#),
      228 => to_slv(opcode_type, 16#10#),
      229 => to_slv(opcode_type, 16#0F#),
      230 => to_slv(opcode_type, 16#06#),
      231 => to_slv(opcode_type, 16#03#),
      232 => to_slv(opcode_type, 16#11#),
      233 => to_slv(opcode_type, 16#02#),
      234 => to_slv(opcode_type, 16#0B#),
      235 => to_slv(opcode_type, 16#08#),
      236 => to_slv(opcode_type, 16#06#),
      237 => to_slv(opcode_type, 16#02#),
      238 => to_slv(opcode_type, 16#10#),
      239 => to_slv(opcode_type, 16#09#),
      240 => to_slv(opcode_type, 16#0A#),
      241 => to_slv(opcode_type, 16#0C#),
      242 => to_slv(opcode_type, 16#07#),
      243 => to_slv(opcode_type, 16#09#),
      244 => to_slv(opcode_type, 16#0D#),
      245 => to_slv(opcode_type, 16#0E#),
      246 => to_slv(opcode_type, 16#08#),
      247 => to_slv(opcode_type, 16#0F#),
      248 => to_slv(opcode_type, 16#0F#),
      249 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#06#),
      257 => to_slv(opcode_type, 16#06#),
      258 => to_slv(opcode_type, 16#03#),
      259 => to_slv(opcode_type, 16#05#),
      260 => to_slv(opcode_type, 16#0D#),
      261 => to_slv(opcode_type, 16#09#),
      262 => to_slv(opcode_type, 16#02#),
      263 => to_slv(opcode_type, 16#10#),
      264 => to_slv(opcode_type, 16#07#),
      265 => to_slv(opcode_type, 16#0F#),
      266 => to_slv(opcode_type, 16#0E#),
      267 => to_slv(opcode_type, 16#08#),
      268 => to_slv(opcode_type, 16#08#),
      269 => to_slv(opcode_type, 16#08#),
      270 => to_slv(opcode_type, 16#11#),
      271 => to_slv(opcode_type, 16#0D#),
      272 => to_slv(opcode_type, 16#07#),
      273 => to_slv(opcode_type, 16#10#),
      274 => to_slv(opcode_type, 16#0A#),
      275 => to_slv(opcode_type, 16#08#),
      276 => to_slv(opcode_type, 16#09#),
      277 => to_slv(opcode_type, 16#0B#),
      278 => to_slv(opcode_type, 16#11#),
      279 => to_slv(opcode_type, 16#04#),
      280 => to_slv(opcode_type, 16#0F#),
      281 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#08#),
      290 => to_slv(opcode_type, 16#05#),
      291 => to_slv(opcode_type, 16#09#),
      292 => to_slv(opcode_type, 16#C6#),
      293 => to_slv(opcode_type, 16#0D#),
      294 => to_slv(opcode_type, 16#01#),
      295 => to_slv(opcode_type, 16#09#),
      296 => to_slv(opcode_type, 16#10#),
      297 => to_slv(opcode_type, 16#0D#),
      298 => to_slv(opcode_type, 16#08#),
      299 => to_slv(opcode_type, 16#07#),
      300 => to_slv(opcode_type, 16#08#),
      301 => to_slv(opcode_type, 16#11#),
      302 => to_slv(opcode_type, 16#10#),
      303 => to_slv(opcode_type, 16#07#),
      304 => to_slv(opcode_type, 16#11#),
      305 => to_slv(opcode_type, 16#8F#),
      306 => to_slv(opcode_type, 16#07#),
      307 => to_slv(opcode_type, 16#07#),
      308 => to_slv(opcode_type, 16#10#),
      309 => to_slv(opcode_type, 16#0F#),
      310 => to_slv(opcode_type, 16#09#),
      311 => to_slv(opcode_type, 16#0E#),
      312 => to_slv(opcode_type, 16#11#),
      313 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#07#),
      321 => to_slv(opcode_type, 16#08#),
      322 => to_slv(opcode_type, 16#01#),
      323 => to_slv(opcode_type, 16#02#),
      324 => to_slv(opcode_type, 16#47#),
      325 => to_slv(opcode_type, 16#08#),
      326 => to_slv(opcode_type, 16#08#),
      327 => to_slv(opcode_type, 16#11#),
      328 => to_slv(opcode_type, 16#0D#),
      329 => to_slv(opcode_type, 16#07#),
      330 => to_slv(opcode_type, 16#0B#),
      331 => to_slv(opcode_type, 16#0E#),
      332 => to_slv(opcode_type, 16#06#),
      333 => to_slv(opcode_type, 16#06#),
      334 => to_slv(opcode_type, 16#09#),
      335 => to_slv(opcode_type, 16#0F#),
      336 => to_slv(opcode_type, 16#0D#),
      337 => to_slv(opcode_type, 16#06#),
      338 => to_slv(opcode_type, 16#0D#),
      339 => to_slv(opcode_type, 16#11#),
      340 => to_slv(opcode_type, 16#09#),
      341 => to_slv(opcode_type, 16#05#),
      342 => to_slv(opcode_type, 16#0A#),
      343 => to_slv(opcode_type, 16#05#),
      344 => to_slv(opcode_type, 16#0E#),
      345 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#06#),
      353 => to_slv(opcode_type, 16#08#),
      354 => to_slv(opcode_type, 16#05#),
      355 => to_slv(opcode_type, 16#03#),
      356 => to_slv(opcode_type, 16#0D#),
      357 => to_slv(opcode_type, 16#09#),
      358 => to_slv(opcode_type, 16#02#),
      359 => to_slv(opcode_type, 16#0B#),
      360 => to_slv(opcode_type, 16#01#),
      361 => to_slv(opcode_type, 16#0B#),
      362 => to_slv(opcode_type, 16#09#),
      363 => to_slv(opcode_type, 16#09#),
      364 => to_slv(opcode_type, 16#08#),
      365 => to_slv(opcode_type, 16#0E#),
      366 => to_slv(opcode_type, 16#0C#),
      367 => to_slv(opcode_type, 16#09#),
      368 => to_slv(opcode_type, 16#11#),
      369 => to_slv(opcode_type, 16#0B#),
      370 => to_slv(opcode_type, 16#07#),
      371 => to_slv(opcode_type, 16#08#),
      372 => to_slv(opcode_type, 16#0F#),
      373 => to_slv(opcode_type, 16#10#),
      374 => to_slv(opcode_type, 16#06#),
      375 => to_slv(opcode_type, 16#0C#),
      376 => to_slv(opcode_type, 16#C9#),
      377 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#06#),
      385 => to_slv(opcode_type, 16#09#),
      386 => to_slv(opcode_type, 16#04#),
      387 => to_slv(opcode_type, 16#03#),
      388 => to_slv(opcode_type, 16#0B#),
      389 => to_slv(opcode_type, 16#06#),
      390 => to_slv(opcode_type, 16#02#),
      391 => to_slv(opcode_type, 16#0E#),
      392 => to_slv(opcode_type, 16#07#),
      393 => to_slv(opcode_type, 16#0F#),
      394 => to_slv(opcode_type, 16#0D#),
      395 => to_slv(opcode_type, 16#09#),
      396 => to_slv(opcode_type, 16#06#),
      397 => to_slv(opcode_type, 16#02#),
      398 => to_slv(opcode_type, 16#0C#),
      399 => to_slv(opcode_type, 16#07#),
      400 => to_slv(opcode_type, 16#3F#),
      401 => to_slv(opcode_type, 16#0A#),
      402 => to_slv(opcode_type, 16#09#),
      403 => to_slv(opcode_type, 16#06#),
      404 => to_slv(opcode_type, 16#11#),
      405 => to_slv(opcode_type, 16#10#),
      406 => to_slv(opcode_type, 16#07#),
      407 => to_slv(opcode_type, 16#0C#),
      408 => to_slv(opcode_type, 16#10#),
      409 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#06#),
      417 => to_slv(opcode_type, 16#08#),
      418 => to_slv(opcode_type, 16#09#),
      419 => to_slv(opcode_type, 16#05#),
      420 => to_slv(opcode_type, 16#0A#),
      421 => to_slv(opcode_type, 16#05#),
      422 => to_slv(opcode_type, 16#0F#),
      423 => to_slv(opcode_type, 16#01#),
      424 => to_slv(opcode_type, 16#03#),
      425 => to_slv(opcode_type, 16#0B#),
      426 => to_slv(opcode_type, 16#07#),
      427 => to_slv(opcode_type, 16#07#),
      428 => to_slv(opcode_type, 16#08#),
      429 => to_slv(opcode_type, 16#11#),
      430 => to_slv(opcode_type, 16#0A#),
      431 => to_slv(opcode_type, 16#07#),
      432 => to_slv(opcode_type, 16#11#),
      433 => to_slv(opcode_type, 16#11#),
      434 => to_slv(opcode_type, 16#07#),
      435 => to_slv(opcode_type, 16#08#),
      436 => to_slv(opcode_type, 16#0C#),
      437 => to_slv(opcode_type, 16#12#),
      438 => to_slv(opcode_type, 16#06#),
      439 => to_slv(opcode_type, 16#0E#),
      440 => to_slv(opcode_type, 16#0C#),
      441 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#07#),
      449 => to_slv(opcode_type, 16#09#),
      450 => to_slv(opcode_type, 16#03#),
      451 => to_slv(opcode_type, 16#02#),
      452 => to_slv(opcode_type, 16#0E#),
      453 => to_slv(opcode_type, 16#09#),
      454 => to_slv(opcode_type, 16#04#),
      455 => to_slv(opcode_type, 16#0D#),
      456 => to_slv(opcode_type, 16#05#),
      457 => to_slv(opcode_type, 16#11#),
      458 => to_slv(opcode_type, 16#06#),
      459 => to_slv(opcode_type, 16#08#),
      460 => to_slv(opcode_type, 16#08#),
      461 => to_slv(opcode_type, 16#10#),
      462 => to_slv(opcode_type, 16#D3#),
      463 => to_slv(opcode_type, 16#07#),
      464 => to_slv(opcode_type, 16#0E#),
      465 => to_slv(opcode_type, 16#0E#),
      466 => to_slv(opcode_type, 16#06#),
      467 => to_slv(opcode_type, 16#07#),
      468 => to_slv(opcode_type, 16#5E#),
      469 => to_slv(opcode_type, 16#B2#),
      470 => to_slv(opcode_type, 16#07#),
      471 => to_slv(opcode_type, 16#A6#),
      472 => to_slv(opcode_type, 16#0E#),
      473 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#08#),
      481 => to_slv(opcode_type, 16#07#),
      482 => to_slv(opcode_type, 16#01#),
      483 => to_slv(opcode_type, 16#06#),
      484 => to_slv(opcode_type, 16#0A#),
      485 => to_slv(opcode_type, 16#10#),
      486 => to_slv(opcode_type, 16#07#),
      487 => to_slv(opcode_type, 16#04#),
      488 => to_slv(opcode_type, 16#0E#),
      489 => to_slv(opcode_type, 16#08#),
      490 => to_slv(opcode_type, 16#0E#),
      491 => to_slv(opcode_type, 16#0F#),
      492 => to_slv(opcode_type, 16#08#),
      493 => to_slv(opcode_type, 16#06#),
      494 => to_slv(opcode_type, 16#04#),
      495 => to_slv(opcode_type, 16#0D#),
      496 => to_slv(opcode_type, 16#02#),
      497 => to_slv(opcode_type, 16#0B#),
      498 => to_slv(opcode_type, 16#08#),
      499 => to_slv(opcode_type, 16#06#),
      500 => to_slv(opcode_type, 16#0B#),
      501 => to_slv(opcode_type, 16#0A#),
      502 => to_slv(opcode_type, 16#08#),
      503 => to_slv(opcode_type, 16#10#),
      504 => to_slv(opcode_type, 16#11#),
      505 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#07#),
      514 => to_slv(opcode_type, 16#08#),
      515 => to_slv(opcode_type, 16#06#),
      516 => to_slv(opcode_type, 16#0F#),
      517 => to_slv(opcode_type, 16#0F#),
      518 => to_slv(opcode_type, 16#06#),
      519 => to_slv(opcode_type, 16#10#),
      520 => to_slv(opcode_type, 16#0D#),
      521 => to_slv(opcode_type, 16#04#),
      522 => to_slv(opcode_type, 16#03#),
      523 => to_slv(opcode_type, 16#0A#),
      524 => to_slv(opcode_type, 16#07#),
      525 => to_slv(opcode_type, 16#08#),
      526 => to_slv(opcode_type, 16#05#),
      527 => to_slv(opcode_type, 16#0B#),
      528 => to_slv(opcode_type, 16#09#),
      529 => to_slv(opcode_type, 16#11#),
      530 => to_slv(opcode_type, 16#42#),
      531 => to_slv(opcode_type, 16#08#),
      532 => to_slv(opcode_type, 16#05#),
      533 => to_slv(opcode_type, 16#0F#),
      534 => to_slv(opcode_type, 16#09#),
      535 => to_slv(opcode_type, 16#0C#),
      536 => to_slv(opcode_type, 16#0E#),
      537 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#09#),
      545 => to_slv(opcode_type, 16#06#),
      546 => to_slv(opcode_type, 16#06#),
      547 => to_slv(opcode_type, 16#08#),
      548 => to_slv(opcode_type, 16#0E#),
      549 => to_slv(opcode_type, 16#11#),
      550 => to_slv(opcode_type, 16#03#),
      551 => to_slv(opcode_type, 16#11#),
      552 => to_slv(opcode_type, 16#08#),
      553 => to_slv(opcode_type, 16#04#),
      554 => to_slv(opcode_type, 16#0A#),
      555 => to_slv(opcode_type, 16#06#),
      556 => to_slv(opcode_type, 16#11#),
      557 => to_slv(opcode_type, 16#0D#),
      558 => to_slv(opcode_type, 16#06#),
      559 => to_slv(opcode_type, 16#04#),
      560 => to_slv(opcode_type, 16#08#),
      561 => to_slv(opcode_type, 16#0A#),
      562 => to_slv(opcode_type, 16#0F#),
      563 => to_slv(opcode_type, 16#06#),
      564 => to_slv(opcode_type, 16#02#),
      565 => to_slv(opcode_type, 16#0B#),
      566 => to_slv(opcode_type, 16#09#),
      567 => to_slv(opcode_type, 16#0D#),
      568 => to_slv(opcode_type, 16#0E#),
      569 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#09#),
      577 => to_slv(opcode_type, 16#08#),
      578 => to_slv(opcode_type, 16#01#),
      579 => to_slv(opcode_type, 16#09#),
      580 => to_slv(opcode_type, 16#11#),
      581 => to_slv(opcode_type, 16#0F#),
      582 => to_slv(opcode_type, 16#07#),
      583 => to_slv(opcode_type, 16#03#),
      584 => to_slv(opcode_type, 16#0C#),
      585 => to_slv(opcode_type, 16#04#),
      586 => to_slv(opcode_type, 16#0C#),
      587 => to_slv(opcode_type, 16#06#),
      588 => to_slv(opcode_type, 16#06#),
      589 => to_slv(opcode_type, 16#02#),
      590 => to_slv(opcode_type, 16#0F#),
      591 => to_slv(opcode_type, 16#07#),
      592 => to_slv(opcode_type, 16#0E#),
      593 => to_slv(opcode_type, 16#49#),
      594 => to_slv(opcode_type, 16#09#),
      595 => to_slv(opcode_type, 16#06#),
      596 => to_slv(opcode_type, 16#0B#),
      597 => to_slv(opcode_type, 16#0A#),
      598 => to_slv(opcode_type, 16#09#),
      599 => to_slv(opcode_type, 16#0E#),
      600 => to_slv(opcode_type, 16#0D#),
      601 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#06#),
      609 => to_slv(opcode_type, 16#08#),
      610 => to_slv(opcode_type, 16#09#),
      611 => to_slv(opcode_type, 16#02#),
      612 => to_slv(opcode_type, 16#0B#),
      613 => to_slv(opcode_type, 16#04#),
      614 => to_slv(opcode_type, 16#11#),
      615 => to_slv(opcode_type, 16#02#),
      616 => to_slv(opcode_type, 16#03#),
      617 => to_slv(opcode_type, 16#0E#),
      618 => to_slv(opcode_type, 16#09#),
      619 => to_slv(opcode_type, 16#08#),
      620 => to_slv(opcode_type, 16#08#),
      621 => to_slv(opcode_type, 16#0A#),
      622 => to_slv(opcode_type, 16#0D#),
      623 => to_slv(opcode_type, 16#07#),
      624 => to_slv(opcode_type, 16#0B#),
      625 => to_slv(opcode_type, 16#0F#),
      626 => to_slv(opcode_type, 16#07#),
      627 => to_slv(opcode_type, 16#08#),
      628 => to_slv(opcode_type, 16#0E#),
      629 => to_slv(opcode_type, 16#0B#),
      630 => to_slv(opcode_type, 16#07#),
      631 => to_slv(opcode_type, 16#0F#),
      632 => to_slv(opcode_type, 16#11#),
      633 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#08#),
      641 => to_slv(opcode_type, 16#07#),
      642 => to_slv(opcode_type, 16#08#),
      643 => to_slv(opcode_type, 16#07#),
      644 => to_slv(opcode_type, 16#10#),
      645 => to_slv(opcode_type, 16#0B#),
      646 => to_slv(opcode_type, 16#02#),
      647 => to_slv(opcode_type, 16#0B#),
      648 => to_slv(opcode_type, 16#07#),
      649 => to_slv(opcode_type, 16#08#),
      650 => to_slv(opcode_type, 16#0E#),
      651 => to_slv(opcode_type, 16#0F#),
      652 => to_slv(opcode_type, 16#05#),
      653 => to_slv(opcode_type, 16#0D#),
      654 => to_slv(opcode_type, 16#06#),
      655 => to_slv(opcode_type, 16#08#),
      656 => to_slv(opcode_type, 16#04#),
      657 => to_slv(opcode_type, 16#0B#),
      658 => to_slv(opcode_type, 16#01#),
      659 => to_slv(opcode_type, 16#0F#),
      660 => to_slv(opcode_type, 16#06#),
      661 => to_slv(opcode_type, 16#02#),
      662 => to_slv(opcode_type, 16#F1#),
      663 => to_slv(opcode_type, 16#01#),
      664 => to_slv(opcode_type, 16#D7#),
      665 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#06#),
      673 => to_slv(opcode_type, 16#09#),
      674 => to_slv(opcode_type, 16#03#),
      675 => to_slv(opcode_type, 16#03#),
      676 => to_slv(opcode_type, 16#13#),
      677 => to_slv(opcode_type, 16#09#),
      678 => to_slv(opcode_type, 16#05#),
      679 => to_slv(opcode_type, 16#0F#),
      680 => to_slv(opcode_type, 16#08#),
      681 => to_slv(opcode_type, 16#0A#),
      682 => to_slv(opcode_type, 16#0A#),
      683 => to_slv(opcode_type, 16#08#),
      684 => to_slv(opcode_type, 16#07#),
      685 => to_slv(opcode_type, 16#04#),
      686 => to_slv(opcode_type, 16#0C#),
      687 => to_slv(opcode_type, 16#07#),
      688 => to_slv(opcode_type, 16#3B#),
      689 => to_slv(opcode_type, 16#0E#),
      690 => to_slv(opcode_type, 16#06#),
      691 => to_slv(opcode_type, 16#07#),
      692 => to_slv(opcode_type, 16#0E#),
      693 => to_slv(opcode_type, 16#0D#),
      694 => to_slv(opcode_type, 16#07#),
      695 => to_slv(opcode_type, 16#0D#),
      696 => to_slv(opcode_type, 16#0D#),
      697 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#07#),
      705 => to_slv(opcode_type, 16#07#),
      706 => to_slv(opcode_type, 16#02#),
      707 => to_slv(opcode_type, 16#07#),
      708 => to_slv(opcode_type, 16#0A#),
      709 => to_slv(opcode_type, 16#0C#),
      710 => to_slv(opcode_type, 16#09#),
      711 => to_slv(opcode_type, 16#02#),
      712 => to_slv(opcode_type, 16#10#),
      713 => to_slv(opcode_type, 16#03#),
      714 => to_slv(opcode_type, 16#0E#),
      715 => to_slv(opcode_type, 16#07#),
      716 => to_slv(opcode_type, 16#09#),
      717 => to_slv(opcode_type, 16#09#),
      718 => to_slv(opcode_type, 16#11#),
      719 => to_slv(opcode_type, 16#0B#),
      720 => to_slv(opcode_type, 16#03#),
      721 => to_slv(opcode_type, 16#0D#),
      722 => to_slv(opcode_type, 16#09#),
      723 => to_slv(opcode_type, 16#09#),
      724 => to_slv(opcode_type, 16#0B#),
      725 => to_slv(opcode_type, 16#11#),
      726 => to_slv(opcode_type, 16#07#),
      727 => to_slv(opcode_type, 16#11#),
      728 => to_slv(opcode_type, 16#0F#),
      729 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#09#),
      737 => to_slv(opcode_type, 16#06#),
      738 => to_slv(opcode_type, 16#08#),
      739 => to_slv(opcode_type, 16#02#),
      740 => to_slv(opcode_type, 16#0C#),
      741 => to_slv(opcode_type, 16#07#),
      742 => to_slv(opcode_type, 16#0C#),
      743 => to_slv(opcode_type, 16#0E#),
      744 => to_slv(opcode_type, 16#08#),
      745 => to_slv(opcode_type, 16#04#),
      746 => to_slv(opcode_type, 16#11#),
      747 => to_slv(opcode_type, 16#06#),
      748 => to_slv(opcode_type, 16#0C#),
      749 => to_slv(opcode_type, 16#0F#),
      750 => to_slv(opcode_type, 16#06#),
      751 => to_slv(opcode_type, 16#01#),
      752 => to_slv(opcode_type, 16#04#),
      753 => to_slv(opcode_type, 16#0C#),
      754 => to_slv(opcode_type, 16#07#),
      755 => to_slv(opcode_type, 16#08#),
      756 => to_slv(opcode_type, 16#0F#),
      757 => to_slv(opcode_type, 16#0D#),
      758 => to_slv(opcode_type, 16#07#),
      759 => to_slv(opcode_type, 16#0E#),
      760 => to_slv(opcode_type, 16#0F#),
      761 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#07#),
      769 => to_slv(opcode_type, 16#06#),
      770 => to_slv(opcode_type, 16#07#),
      771 => to_slv(opcode_type, 16#08#),
      772 => to_slv(opcode_type, 16#0B#),
      773 => to_slv(opcode_type, 16#0A#),
      774 => to_slv(opcode_type, 16#04#),
      775 => to_slv(opcode_type, 16#0B#),
      776 => to_slv(opcode_type, 16#04#),
      777 => to_slv(opcode_type, 16#02#),
      778 => to_slv(opcode_type, 16#0E#),
      779 => to_slv(opcode_type, 16#06#),
      780 => to_slv(opcode_type, 16#06#),
      781 => to_slv(opcode_type, 16#06#),
      782 => to_slv(opcode_type, 16#10#),
      783 => to_slv(opcode_type, 16#0B#),
      784 => to_slv(opcode_type, 16#09#),
      785 => to_slv(opcode_type, 16#10#),
      786 => to_slv(opcode_type, 16#2E#),
      787 => to_slv(opcode_type, 16#08#),
      788 => to_slv(opcode_type, 16#03#),
      789 => to_slv(opcode_type, 16#91#),
      790 => to_slv(opcode_type, 16#06#),
      791 => to_slv(opcode_type, 16#10#),
      792 => to_slv(opcode_type, 16#0F#),
      793 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#08#),
      801 => to_slv(opcode_type, 16#08#),
      802 => to_slv(opcode_type, 16#04#),
      803 => to_slv(opcode_type, 16#08#),
      804 => to_slv(opcode_type, 16#0D#),
      805 => to_slv(opcode_type, 16#0A#),
      806 => to_slv(opcode_type, 16#08#),
      807 => to_slv(opcode_type, 16#01#),
      808 => to_slv(opcode_type, 16#0A#),
      809 => to_slv(opcode_type, 16#09#),
      810 => to_slv(opcode_type, 16#0B#),
      811 => to_slv(opcode_type, 16#0D#),
      812 => to_slv(opcode_type, 16#07#),
      813 => to_slv(opcode_type, 16#06#),
      814 => to_slv(opcode_type, 16#09#),
      815 => to_slv(opcode_type, 16#0C#),
      816 => to_slv(opcode_type, 16#10#),
      817 => to_slv(opcode_type, 16#05#),
      818 => to_slv(opcode_type, 16#10#),
      819 => to_slv(opcode_type, 16#06#),
      820 => to_slv(opcode_type, 16#07#),
      821 => to_slv(opcode_type, 16#11#),
      822 => to_slv(opcode_type, 16#10#),
      823 => to_slv(opcode_type, 16#01#),
      824 => to_slv(opcode_type, 16#0D#),
      825 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#07#),
      833 => to_slv(opcode_type, 16#06#),
      834 => to_slv(opcode_type, 16#09#),
      835 => to_slv(opcode_type, 16#09#),
      836 => to_slv(opcode_type, 16#0C#),
      837 => to_slv(opcode_type, 16#C6#),
      838 => to_slv(opcode_type, 16#06#),
      839 => to_slv(opcode_type, 16#10#),
      840 => to_slv(opcode_type, 16#0A#),
      841 => to_slv(opcode_type, 16#02#),
      842 => to_slv(opcode_type, 16#09#),
      843 => to_slv(opcode_type, 16#0E#),
      844 => to_slv(opcode_type, 16#FD#),
      845 => to_slv(opcode_type, 16#09#),
      846 => to_slv(opcode_type, 16#01#),
      847 => to_slv(opcode_type, 16#06#),
      848 => to_slv(opcode_type, 16#10#),
      849 => to_slv(opcode_type, 16#0C#),
      850 => to_slv(opcode_type, 16#06#),
      851 => to_slv(opcode_type, 16#06#),
      852 => to_slv(opcode_type, 16#0B#),
      853 => to_slv(opcode_type, 16#0A#),
      854 => to_slv(opcode_type, 16#09#),
      855 => to_slv(opcode_type, 16#10#),
      856 => to_slv(opcode_type, 16#0B#),
      857 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#09#),
      865 => to_slv(opcode_type, 16#07#),
      866 => to_slv(opcode_type, 16#07#),
      867 => to_slv(opcode_type, 16#07#),
      868 => to_slv(opcode_type, 16#0A#),
      869 => to_slv(opcode_type, 16#0D#),
      870 => to_slv(opcode_type, 16#09#),
      871 => to_slv(opcode_type, 16#0E#),
      872 => to_slv(opcode_type, 16#0A#),
      873 => to_slv(opcode_type, 16#02#),
      874 => to_slv(opcode_type, 16#01#),
      875 => to_slv(opcode_type, 16#0C#),
      876 => to_slv(opcode_type, 16#07#),
      877 => to_slv(opcode_type, 16#07#),
      878 => to_slv(opcode_type, 16#07#),
      879 => to_slv(opcode_type, 16#0F#),
      880 => to_slv(opcode_type, 16#0B#),
      881 => to_slv(opcode_type, 16#07#),
      882 => to_slv(opcode_type, 16#11#),
      883 => to_slv(opcode_type, 16#C5#),
      884 => to_slv(opcode_type, 16#09#),
      885 => to_slv(opcode_type, 16#06#),
      886 => to_slv(opcode_type, 16#0F#),
      887 => to_slv(opcode_type, 16#0C#),
      888 => to_slv(opcode_type, 16#11#),
      889 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#08#),
      897 => to_slv(opcode_type, 16#09#),
      898 => to_slv(opcode_type, 16#09#),
      899 => to_slv(opcode_type, 16#01#),
      900 => to_slv(opcode_type, 16#0D#),
      901 => to_slv(opcode_type, 16#01#),
      902 => to_slv(opcode_type, 16#0B#),
      903 => to_slv(opcode_type, 16#01#),
      904 => to_slv(opcode_type, 16#05#),
      905 => to_slv(opcode_type, 16#10#),
      906 => to_slv(opcode_type, 16#08#),
      907 => to_slv(opcode_type, 16#09#),
      908 => to_slv(opcode_type, 16#07#),
      909 => to_slv(opcode_type, 16#4B#),
      910 => to_slv(opcode_type, 16#0A#),
      911 => to_slv(opcode_type, 16#09#),
      912 => to_slv(opcode_type, 16#0D#),
      913 => to_slv(opcode_type, 16#0B#),
      914 => to_slv(opcode_type, 16#08#),
      915 => to_slv(opcode_type, 16#07#),
      916 => to_slv(opcode_type, 16#45#),
      917 => to_slv(opcode_type, 16#0E#),
      918 => to_slv(opcode_type, 16#07#),
      919 => to_slv(opcode_type, 16#10#),
      920 => to_slv(opcode_type, 16#0F#),
      921 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#08#),
      929 => to_slv(opcode_type, 16#09#),
      930 => to_slv(opcode_type, 16#09#),
      931 => to_slv(opcode_type, 16#08#),
      932 => to_slv(opcode_type, 16#0A#),
      933 => to_slv(opcode_type, 16#10#),
      934 => to_slv(opcode_type, 16#01#),
      935 => to_slv(opcode_type, 16#0D#),
      936 => to_slv(opcode_type, 16#04#),
      937 => to_slv(opcode_type, 16#07#),
      938 => to_slv(opcode_type, 16#11#),
      939 => to_slv(opcode_type, 16#22#),
      940 => to_slv(opcode_type, 16#07#),
      941 => to_slv(opcode_type, 16#07#),
      942 => to_slv(opcode_type, 16#09#),
      943 => to_slv(opcode_type, 16#10#),
      944 => to_slv(opcode_type, 16#0A#),
      945 => to_slv(opcode_type, 16#08#),
      946 => to_slv(opcode_type, 16#0C#),
      947 => to_slv(opcode_type, 16#0C#),
      948 => to_slv(opcode_type, 16#09#),
      949 => to_slv(opcode_type, 16#07#),
      950 => to_slv(opcode_type, 16#9B#),
      951 => to_slv(opcode_type, 16#0A#),
      952 => to_slv(opcode_type, 16#11#),
      953 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#09#),
      962 => to_slv(opcode_type, 16#01#),
      963 => to_slv(opcode_type, 16#02#),
      964 => to_slv(opcode_type, 16#0C#),
      965 => to_slv(opcode_type, 16#06#),
      966 => to_slv(opcode_type, 16#04#),
      967 => to_slv(opcode_type, 16#10#),
      968 => to_slv(opcode_type, 16#06#),
      969 => to_slv(opcode_type, 16#0A#),
      970 => to_slv(opcode_type, 16#0A#),
      971 => to_slv(opcode_type, 16#09#),
      972 => to_slv(opcode_type, 16#09#),
      973 => to_slv(opcode_type, 16#01#),
      974 => to_slv(opcode_type, 16#0C#),
      975 => to_slv(opcode_type, 16#09#),
      976 => to_slv(opcode_type, 16#C3#),
      977 => to_slv(opcode_type, 16#0E#),
      978 => to_slv(opcode_type, 16#09#),
      979 => to_slv(opcode_type, 16#08#),
      980 => to_slv(opcode_type, 16#0B#),
      981 => to_slv(opcode_type, 16#0A#),
      982 => to_slv(opcode_type, 16#08#),
      983 => to_slv(opcode_type, 16#0A#),
      984 => to_slv(opcode_type, 16#11#),
      985 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#06#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#07#),
      995 => to_slv(opcode_type, 16#05#),
      996 => to_slv(opcode_type, 16#70#),
      997 => to_slv(opcode_type, 16#01#),
      998 => to_slv(opcode_type, 16#E2#),
      999 => to_slv(opcode_type, 16#04#),
      1000 => to_slv(opcode_type, 16#07#),
      1001 => to_slv(opcode_type, 16#0C#),
      1002 => to_slv(opcode_type, 16#0A#),
      1003 => to_slv(opcode_type, 16#07#),
      1004 => to_slv(opcode_type, 16#06#),
      1005 => to_slv(opcode_type, 16#03#),
      1006 => to_slv(opcode_type, 16#0D#),
      1007 => to_slv(opcode_type, 16#07#),
      1008 => to_slv(opcode_type, 16#0E#),
      1009 => to_slv(opcode_type, 16#10#),
      1010 => to_slv(opcode_type, 16#06#),
      1011 => to_slv(opcode_type, 16#08#),
      1012 => to_slv(opcode_type, 16#0D#),
      1013 => to_slv(opcode_type, 16#0B#),
      1014 => to_slv(opcode_type, 16#06#),
      1015 => to_slv(opcode_type, 16#11#),
      1016 => to_slv(opcode_type, 16#51#),
      1017 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#07#),
      1025 => to_slv(opcode_type, 16#07#),
      1026 => to_slv(opcode_type, 16#07#),
      1027 => to_slv(opcode_type, 16#08#),
      1028 => to_slv(opcode_type, 16#0C#),
      1029 => to_slv(opcode_type, 16#0B#),
      1030 => to_slv(opcode_type, 16#06#),
      1031 => to_slv(opcode_type, 16#0E#),
      1032 => to_slv(opcode_type, 16#0C#),
      1033 => to_slv(opcode_type, 16#04#),
      1034 => to_slv(opcode_type, 16#08#),
      1035 => to_slv(opcode_type, 16#0F#),
      1036 => to_slv(opcode_type, 16#0F#),
      1037 => to_slv(opcode_type, 16#08#),
      1038 => to_slv(opcode_type, 16#05#),
      1039 => to_slv(opcode_type, 16#07#),
      1040 => to_slv(opcode_type, 16#0C#),
      1041 => to_slv(opcode_type, 16#0B#),
      1042 => to_slv(opcode_type, 16#08#),
      1043 => to_slv(opcode_type, 16#06#),
      1044 => to_slv(opcode_type, 16#0A#),
      1045 => to_slv(opcode_type, 16#11#),
      1046 => to_slv(opcode_type, 16#07#),
      1047 => to_slv(opcode_type, 16#0E#),
      1048 => to_slv(opcode_type, 16#3C#),
      1049 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#09#),
      1057 => to_slv(opcode_type, 16#07#),
      1058 => to_slv(opcode_type, 16#05#),
      1059 => to_slv(opcode_type, 16#08#),
      1060 => to_slv(opcode_type, 16#0E#),
      1061 => to_slv(opcode_type, 16#10#),
      1062 => to_slv(opcode_type, 16#01#),
      1063 => to_slv(opcode_type, 16#09#),
      1064 => to_slv(opcode_type, 16#0F#),
      1065 => to_slv(opcode_type, 16#0E#),
      1066 => to_slv(opcode_type, 16#06#),
      1067 => to_slv(opcode_type, 16#06#),
      1068 => to_slv(opcode_type, 16#09#),
      1069 => to_slv(opcode_type, 16#0E#),
      1070 => to_slv(opcode_type, 16#0C#),
      1071 => to_slv(opcode_type, 16#09#),
      1072 => to_slv(opcode_type, 16#10#),
      1073 => to_slv(opcode_type, 16#0C#),
      1074 => to_slv(opcode_type, 16#09#),
      1075 => to_slv(opcode_type, 16#09#),
      1076 => to_slv(opcode_type, 16#0E#),
      1077 => to_slv(opcode_type, 16#0A#),
      1078 => to_slv(opcode_type, 16#08#),
      1079 => to_slv(opcode_type, 16#0E#),
      1080 => to_slv(opcode_type, 16#11#),
      1081 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#08#),
      1089 => to_slv(opcode_type, 16#06#),
      1090 => to_slv(opcode_type, 16#04#),
      1091 => to_slv(opcode_type, 16#03#),
      1092 => to_slv(opcode_type, 16#0B#),
      1093 => to_slv(opcode_type, 16#08#),
      1094 => to_slv(opcode_type, 16#08#),
      1095 => to_slv(opcode_type, 16#10#),
      1096 => to_slv(opcode_type, 16#0B#),
      1097 => to_slv(opcode_type, 16#03#),
      1098 => to_slv(opcode_type, 16#DB#),
      1099 => to_slv(opcode_type, 16#07#),
      1100 => to_slv(opcode_type, 16#07#),
      1101 => to_slv(opcode_type, 16#03#),
      1102 => to_slv(opcode_type, 16#0D#),
      1103 => to_slv(opcode_type, 16#09#),
      1104 => to_slv(opcode_type, 16#0D#),
      1105 => to_slv(opcode_type, 16#0A#),
      1106 => to_slv(opcode_type, 16#09#),
      1107 => to_slv(opcode_type, 16#06#),
      1108 => to_slv(opcode_type, 16#0A#),
      1109 => to_slv(opcode_type, 16#0B#),
      1110 => to_slv(opcode_type, 16#07#),
      1111 => to_slv(opcode_type, 16#5F#),
      1112 => to_slv(opcode_type, 16#0C#),
      1113 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#09#),
      1121 => to_slv(opcode_type, 16#09#),
      1122 => to_slv(opcode_type, 16#06#),
      1123 => to_slv(opcode_type, 16#08#),
      1124 => to_slv(opcode_type, 16#0D#),
      1125 => to_slv(opcode_type, 16#10#),
      1126 => to_slv(opcode_type, 16#09#),
      1127 => to_slv(opcode_type, 16#0B#),
      1128 => to_slv(opcode_type, 16#0A#),
      1129 => to_slv(opcode_type, 16#01#),
      1130 => to_slv(opcode_type, 16#08#),
      1131 => to_slv(opcode_type, 16#0E#),
      1132 => to_slv(opcode_type, 16#0A#),
      1133 => to_slv(opcode_type, 16#08#),
      1134 => to_slv(opcode_type, 16#05#),
      1135 => to_slv(opcode_type, 16#08#),
      1136 => to_slv(opcode_type, 16#0B#),
      1137 => to_slv(opcode_type, 16#0E#),
      1138 => to_slv(opcode_type, 16#09#),
      1139 => to_slv(opcode_type, 16#07#),
      1140 => to_slv(opcode_type, 16#15#),
      1141 => to_slv(opcode_type, 16#11#),
      1142 => to_slv(opcode_type, 16#08#),
      1143 => to_slv(opcode_type, 16#0A#),
      1144 => to_slv(opcode_type, 16#0D#),
      1145 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#08#),
      1153 => to_slv(opcode_type, 16#09#),
      1154 => to_slv(opcode_type, 16#02#),
      1155 => to_slv(opcode_type, 16#07#),
      1156 => to_slv(opcode_type, 16#11#),
      1157 => to_slv(opcode_type, 16#0C#),
      1158 => to_slv(opcode_type, 16#06#),
      1159 => to_slv(opcode_type, 16#03#),
      1160 => to_slv(opcode_type, 16#0C#),
      1161 => to_slv(opcode_type, 16#04#),
      1162 => to_slv(opcode_type, 16#0A#),
      1163 => to_slv(opcode_type, 16#07#),
      1164 => to_slv(opcode_type, 16#09#),
      1165 => to_slv(opcode_type, 16#05#),
      1166 => to_slv(opcode_type, 16#0E#),
      1167 => to_slv(opcode_type, 16#09#),
      1168 => to_slv(opcode_type, 16#0F#),
      1169 => to_slv(opcode_type, 16#0A#),
      1170 => to_slv(opcode_type, 16#08#),
      1171 => to_slv(opcode_type, 16#08#),
      1172 => to_slv(opcode_type, 16#10#),
      1173 => to_slv(opcode_type, 16#0E#),
      1174 => to_slv(opcode_type, 16#08#),
      1175 => to_slv(opcode_type, 16#0F#),
      1176 => to_slv(opcode_type, 16#11#),
      1177 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#09#),
      1185 => to_slv(opcode_type, 16#07#),
      1186 => to_slv(opcode_type, 16#07#),
      1187 => to_slv(opcode_type, 16#05#),
      1188 => to_slv(opcode_type, 16#0B#),
      1189 => to_slv(opcode_type, 16#02#),
      1190 => to_slv(opcode_type, 16#0F#),
      1191 => to_slv(opcode_type, 16#01#),
      1192 => to_slv(opcode_type, 16#01#),
      1193 => to_slv(opcode_type, 16#0A#),
      1194 => to_slv(opcode_type, 16#08#),
      1195 => to_slv(opcode_type, 16#07#),
      1196 => to_slv(opcode_type, 16#07#),
      1197 => to_slv(opcode_type, 16#0B#),
      1198 => to_slv(opcode_type, 16#BE#),
      1199 => to_slv(opcode_type, 16#09#),
      1200 => to_slv(opcode_type, 16#0E#),
      1201 => to_slv(opcode_type, 16#0A#),
      1202 => to_slv(opcode_type, 16#06#),
      1203 => to_slv(opcode_type, 16#09#),
      1204 => to_slv(opcode_type, 16#0C#),
      1205 => to_slv(opcode_type, 16#0F#),
      1206 => to_slv(opcode_type, 16#06#),
      1207 => to_slv(opcode_type, 16#0B#),
      1208 => to_slv(opcode_type, 16#0B#),
      1209 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#09#),
      1217 => to_slv(opcode_type, 16#06#),
      1218 => to_slv(opcode_type, 16#09#),
      1219 => to_slv(opcode_type, 16#09#),
      1220 => to_slv(opcode_type, 16#4A#),
      1221 => to_slv(opcode_type, 16#0E#),
      1222 => to_slv(opcode_type, 16#08#),
      1223 => to_slv(opcode_type, 16#0E#),
      1224 => to_slv(opcode_type, 16#1C#),
      1225 => to_slv(opcode_type, 16#06#),
      1226 => to_slv(opcode_type, 16#04#),
      1227 => to_slv(opcode_type, 16#B3#),
      1228 => to_slv(opcode_type, 16#09#),
      1229 => to_slv(opcode_type, 16#0A#),
      1230 => to_slv(opcode_type, 16#11#),
      1231 => to_slv(opcode_type, 16#08#),
      1232 => to_slv(opcode_type, 16#02#),
      1233 => to_slv(opcode_type, 16#09#),
      1234 => to_slv(opcode_type, 16#0D#),
      1235 => to_slv(opcode_type, 16#0D#),
      1236 => to_slv(opcode_type, 16#07#),
      1237 => to_slv(opcode_type, 16#03#),
      1238 => to_slv(opcode_type, 16#11#),
      1239 => to_slv(opcode_type, 16#03#),
      1240 => to_slv(opcode_type, 16#0A#),
      1241 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#09#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#01#),
      1251 => to_slv(opcode_type, 16#08#),
      1252 => to_slv(opcode_type, 16#0D#),
      1253 => to_slv(opcode_type, 16#11#),
      1254 => to_slv(opcode_type, 16#07#),
      1255 => to_slv(opcode_type, 16#08#),
      1256 => to_slv(opcode_type, 16#0D#),
      1257 => to_slv(opcode_type, 16#0F#),
      1258 => to_slv(opcode_type, 16#01#),
      1259 => to_slv(opcode_type, 16#0E#),
      1260 => to_slv(opcode_type, 16#07#),
      1261 => to_slv(opcode_type, 16#06#),
      1262 => to_slv(opcode_type, 16#01#),
      1263 => to_slv(opcode_type, 16#0E#),
      1264 => to_slv(opcode_type, 16#06#),
      1265 => to_slv(opcode_type, 16#0C#),
      1266 => to_slv(opcode_type, 16#0D#),
      1267 => to_slv(opcode_type, 16#07#),
      1268 => to_slv(opcode_type, 16#07#),
      1269 => to_slv(opcode_type, 16#0F#),
      1270 => to_slv(opcode_type, 16#0A#),
      1271 => to_slv(opcode_type, 16#05#),
      1272 => to_slv(opcode_type, 16#52#),
      1273 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#08#),
      1282 => to_slv(opcode_type, 16#02#),
      1283 => to_slv(opcode_type, 16#07#),
      1284 => to_slv(opcode_type, 16#0B#),
      1285 => to_slv(opcode_type, 16#D5#),
      1286 => to_slv(opcode_type, 16#01#),
      1287 => to_slv(opcode_type, 16#09#),
      1288 => to_slv(opcode_type, 16#0A#),
      1289 => to_slv(opcode_type, 16#0D#),
      1290 => to_slv(opcode_type, 16#07#),
      1291 => to_slv(opcode_type, 16#07#),
      1292 => to_slv(opcode_type, 16#06#),
      1293 => to_slv(opcode_type, 16#0D#),
      1294 => to_slv(opcode_type, 16#10#),
      1295 => to_slv(opcode_type, 16#09#),
      1296 => to_slv(opcode_type, 16#0E#),
      1297 => to_slv(opcode_type, 16#0D#),
      1298 => to_slv(opcode_type, 16#06#),
      1299 => to_slv(opcode_type, 16#09#),
      1300 => to_slv(opcode_type, 16#10#),
      1301 => to_slv(opcode_type, 16#10#),
      1302 => to_slv(opcode_type, 16#08#),
      1303 => to_slv(opcode_type, 16#0A#),
      1304 => to_slv(opcode_type, 16#0C#),
      1305 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#09#),
      1313 => to_slv(opcode_type, 16#06#),
      1314 => to_slv(opcode_type, 16#01#),
      1315 => to_slv(opcode_type, 16#02#),
      1316 => to_slv(opcode_type, 16#0F#),
      1317 => to_slv(opcode_type, 16#06#),
      1318 => to_slv(opcode_type, 16#02#),
      1319 => to_slv(opcode_type, 16#0D#),
      1320 => to_slv(opcode_type, 16#05#),
      1321 => to_slv(opcode_type, 16#0F#),
      1322 => to_slv(opcode_type, 16#07#),
      1323 => to_slv(opcode_type, 16#06#),
      1324 => to_slv(opcode_type, 16#07#),
      1325 => to_slv(opcode_type, 16#0C#),
      1326 => to_slv(opcode_type, 16#0D#),
      1327 => to_slv(opcode_type, 16#07#),
      1328 => to_slv(opcode_type, 16#11#),
      1329 => to_slv(opcode_type, 16#0B#),
      1330 => to_slv(opcode_type, 16#06#),
      1331 => to_slv(opcode_type, 16#06#),
      1332 => to_slv(opcode_type, 16#0D#),
      1333 => to_slv(opcode_type, 16#0A#),
      1334 => to_slv(opcode_type, 16#07#),
      1335 => to_slv(opcode_type, 16#0B#),
      1336 => to_slv(opcode_type, 16#35#),
      1337 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#06#),
      1345 => to_slv(opcode_type, 16#07#),
      1346 => to_slv(opcode_type, 16#05#),
      1347 => to_slv(opcode_type, 16#09#),
      1348 => to_slv(opcode_type, 16#0C#),
      1349 => to_slv(opcode_type, 16#0B#),
      1350 => to_slv(opcode_type, 16#03#),
      1351 => to_slv(opcode_type, 16#06#),
      1352 => to_slv(opcode_type, 16#0F#),
      1353 => to_slv(opcode_type, 16#0F#),
      1354 => to_slv(opcode_type, 16#06#),
      1355 => to_slv(opcode_type, 16#06#),
      1356 => to_slv(opcode_type, 16#06#),
      1357 => to_slv(opcode_type, 16#51#),
      1358 => to_slv(opcode_type, 16#11#),
      1359 => to_slv(opcode_type, 16#06#),
      1360 => to_slv(opcode_type, 16#0C#),
      1361 => to_slv(opcode_type, 16#0C#),
      1362 => to_slv(opcode_type, 16#08#),
      1363 => to_slv(opcode_type, 16#07#),
      1364 => to_slv(opcode_type, 16#11#),
      1365 => to_slv(opcode_type, 16#11#),
      1366 => to_slv(opcode_type, 16#09#),
      1367 => to_slv(opcode_type, 16#0B#),
      1368 => to_slv(opcode_type, 16#0E#),
      1369 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#09#),
      1377 => to_slv(opcode_type, 16#08#),
      1378 => to_slv(opcode_type, 16#02#),
      1379 => to_slv(opcode_type, 16#02#),
      1380 => to_slv(opcode_type, 16#10#),
      1381 => to_slv(opcode_type, 16#09#),
      1382 => to_slv(opcode_type, 16#02#),
      1383 => to_slv(opcode_type, 16#0D#),
      1384 => to_slv(opcode_type, 16#05#),
      1385 => to_slv(opcode_type, 16#0A#),
      1386 => to_slv(opcode_type, 16#07#),
      1387 => to_slv(opcode_type, 16#09#),
      1388 => to_slv(opcode_type, 16#08#),
      1389 => to_slv(opcode_type, 16#0C#),
      1390 => to_slv(opcode_type, 16#0A#),
      1391 => to_slv(opcode_type, 16#08#),
      1392 => to_slv(opcode_type, 16#75#),
      1393 => to_slv(opcode_type, 16#0E#),
      1394 => to_slv(opcode_type, 16#06#),
      1395 => to_slv(opcode_type, 16#09#),
      1396 => to_slv(opcode_type, 16#0E#),
      1397 => to_slv(opcode_type, 16#0E#),
      1398 => to_slv(opcode_type, 16#08#),
      1399 => to_slv(opcode_type, 16#0E#),
      1400 => to_slv(opcode_type, 16#0D#),
      1401 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#08#),
      1410 => to_slv(opcode_type, 16#09#),
      1411 => to_slv(opcode_type, 16#03#),
      1412 => to_slv(opcode_type, 16#0D#),
      1413 => to_slv(opcode_type, 16#09#),
      1414 => to_slv(opcode_type, 16#0A#),
      1415 => to_slv(opcode_type, 16#11#),
      1416 => to_slv(opcode_type, 16#07#),
      1417 => to_slv(opcode_type, 16#07#),
      1418 => to_slv(opcode_type, 16#0F#),
      1419 => to_slv(opcode_type, 16#39#),
      1420 => to_slv(opcode_type, 16#06#),
      1421 => to_slv(opcode_type, 16#0F#),
      1422 => to_slv(opcode_type, 16#0F#),
      1423 => to_slv(opcode_type, 16#08#),
      1424 => to_slv(opcode_type, 16#03#),
      1425 => to_slv(opcode_type, 16#03#),
      1426 => to_slv(opcode_type, 16#0B#),
      1427 => to_slv(opcode_type, 16#06#),
      1428 => to_slv(opcode_type, 16#04#),
      1429 => to_slv(opcode_type, 16#F4#),
      1430 => to_slv(opcode_type, 16#06#),
      1431 => to_slv(opcode_type, 16#0B#),
      1432 => to_slv(opcode_type, 16#DD#),
      1433 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#08#),
      1441 => to_slv(opcode_type, 16#09#),
      1442 => to_slv(opcode_type, 16#02#),
      1443 => to_slv(opcode_type, 16#07#),
      1444 => to_slv(opcode_type, 16#11#),
      1445 => to_slv(opcode_type, 16#0D#),
      1446 => to_slv(opcode_type, 16#05#),
      1447 => to_slv(opcode_type, 16#08#),
      1448 => to_slv(opcode_type, 16#0E#),
      1449 => to_slv(opcode_type, 16#0B#),
      1450 => to_slv(opcode_type, 16#09#),
      1451 => to_slv(opcode_type, 16#07#),
      1452 => to_slv(opcode_type, 16#08#),
      1453 => to_slv(opcode_type, 16#0E#),
      1454 => to_slv(opcode_type, 16#11#),
      1455 => to_slv(opcode_type, 16#06#),
      1456 => to_slv(opcode_type, 16#0B#),
      1457 => to_slv(opcode_type, 16#1F#),
      1458 => to_slv(opcode_type, 16#06#),
      1459 => to_slv(opcode_type, 16#06#),
      1460 => to_slv(opcode_type, 16#0F#),
      1461 => to_slv(opcode_type, 16#0C#),
      1462 => to_slv(opcode_type, 16#09#),
      1463 => to_slv(opcode_type, 16#0F#),
      1464 => to_slv(opcode_type, 16#0B#),
      1465 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#07#),
      1473 => to_slv(opcode_type, 16#07#),
      1474 => to_slv(opcode_type, 16#09#),
      1475 => to_slv(opcode_type, 16#03#),
      1476 => to_slv(opcode_type, 16#0C#),
      1477 => to_slv(opcode_type, 16#09#),
      1478 => to_slv(opcode_type, 16#11#),
      1479 => to_slv(opcode_type, 16#0C#),
      1480 => to_slv(opcode_type, 16#04#),
      1481 => to_slv(opcode_type, 16#08#),
      1482 => to_slv(opcode_type, 16#F0#),
      1483 => to_slv(opcode_type, 16#0F#),
      1484 => to_slv(opcode_type, 16#06#),
      1485 => to_slv(opcode_type, 16#09#),
      1486 => to_slv(opcode_type, 16#09#),
      1487 => to_slv(opcode_type, 16#0C#),
      1488 => to_slv(opcode_type, 16#0A#),
      1489 => to_slv(opcode_type, 16#08#),
      1490 => to_slv(opcode_type, 16#0B#),
      1491 => to_slv(opcode_type, 16#0A#),
      1492 => to_slv(opcode_type, 16#06#),
      1493 => to_slv(opcode_type, 16#05#),
      1494 => to_slv(opcode_type, 16#0E#),
      1495 => to_slv(opcode_type, 16#05#),
      1496 => to_slv(opcode_type, 16#0C#),
      1497 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#07#),
      1505 => to_slv(opcode_type, 16#09#),
      1506 => to_slv(opcode_type, 16#02#),
      1507 => to_slv(opcode_type, 16#04#),
      1508 => to_slv(opcode_type, 16#0C#),
      1509 => to_slv(opcode_type, 16#08#),
      1510 => to_slv(opcode_type, 16#05#),
      1511 => to_slv(opcode_type, 16#0F#),
      1512 => to_slv(opcode_type, 16#05#),
      1513 => to_slv(opcode_type, 16#0E#),
      1514 => to_slv(opcode_type, 16#07#),
      1515 => to_slv(opcode_type, 16#07#),
      1516 => to_slv(opcode_type, 16#09#),
      1517 => to_slv(opcode_type, 16#0B#),
      1518 => to_slv(opcode_type, 16#0C#),
      1519 => to_slv(opcode_type, 16#06#),
      1520 => to_slv(opcode_type, 16#11#),
      1521 => to_slv(opcode_type, 16#0F#),
      1522 => to_slv(opcode_type, 16#08#),
      1523 => to_slv(opcode_type, 16#09#),
      1524 => to_slv(opcode_type, 16#0D#),
      1525 => to_slv(opcode_type, 16#0A#),
      1526 => to_slv(opcode_type, 16#07#),
      1527 => to_slv(opcode_type, 16#0B#),
      1528 => to_slv(opcode_type, 16#0A#),
      1529 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#07#),
      1537 => to_slv(opcode_type, 16#07#),
      1538 => to_slv(opcode_type, 16#04#),
      1539 => to_slv(opcode_type, 16#02#),
      1540 => to_slv(opcode_type, 16#0E#),
      1541 => to_slv(opcode_type, 16#06#),
      1542 => to_slv(opcode_type, 16#04#),
      1543 => to_slv(opcode_type, 16#0F#),
      1544 => to_slv(opcode_type, 16#05#),
      1545 => to_slv(opcode_type, 16#0D#),
      1546 => to_slv(opcode_type, 16#08#),
      1547 => to_slv(opcode_type, 16#09#),
      1548 => to_slv(opcode_type, 16#07#),
      1549 => to_slv(opcode_type, 16#0E#),
      1550 => to_slv(opcode_type, 16#11#),
      1551 => to_slv(opcode_type, 16#07#),
      1552 => to_slv(opcode_type, 16#0A#),
      1553 => to_slv(opcode_type, 16#0A#),
      1554 => to_slv(opcode_type, 16#07#),
      1555 => to_slv(opcode_type, 16#09#),
      1556 => to_slv(opcode_type, 16#0E#),
      1557 => to_slv(opcode_type, 16#CE#),
      1558 => to_slv(opcode_type, 16#08#),
      1559 => to_slv(opcode_type, 16#0E#),
      1560 => to_slv(opcode_type, 16#B4#),
      1561 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#06#),
      1569 => to_slv(opcode_type, 16#07#),
      1570 => to_slv(opcode_type, 16#09#),
      1571 => to_slv(opcode_type, 16#09#),
      1572 => to_slv(opcode_type, 16#11#),
      1573 => to_slv(opcode_type, 16#0F#),
      1574 => to_slv(opcode_type, 16#01#),
      1575 => to_slv(opcode_type, 16#F6#),
      1576 => to_slv(opcode_type, 16#05#),
      1577 => to_slv(opcode_type, 16#08#),
      1578 => to_slv(opcode_type, 16#0A#),
      1579 => to_slv(opcode_type, 16#11#),
      1580 => to_slv(opcode_type, 16#08#),
      1581 => to_slv(opcode_type, 16#09#),
      1582 => to_slv(opcode_type, 16#04#),
      1583 => to_slv(opcode_type, 16#11#),
      1584 => to_slv(opcode_type, 16#04#),
      1585 => to_slv(opcode_type, 16#10#),
      1586 => to_slv(opcode_type, 16#07#),
      1587 => to_slv(opcode_type, 16#07#),
      1588 => to_slv(opcode_type, 16#10#),
      1589 => to_slv(opcode_type, 16#11#),
      1590 => to_slv(opcode_type, 16#09#),
      1591 => to_slv(opcode_type, 16#0F#),
      1592 => to_slv(opcode_type, 16#0D#),
      1593 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#07#),
      1601 => to_slv(opcode_type, 16#08#),
      1602 => to_slv(opcode_type, 16#05#),
      1603 => to_slv(opcode_type, 16#06#),
      1604 => to_slv(opcode_type, 16#10#),
      1605 => to_slv(opcode_type, 16#0C#),
      1606 => to_slv(opcode_type, 16#05#),
      1607 => to_slv(opcode_type, 16#08#),
      1608 => to_slv(opcode_type, 16#11#),
      1609 => to_slv(opcode_type, 16#0A#),
      1610 => to_slv(opcode_type, 16#08#),
      1611 => to_slv(opcode_type, 16#07#),
      1612 => to_slv(opcode_type, 16#06#),
      1613 => to_slv(opcode_type, 16#10#),
      1614 => to_slv(opcode_type, 16#0C#),
      1615 => to_slv(opcode_type, 16#08#),
      1616 => to_slv(opcode_type, 16#2F#),
      1617 => to_slv(opcode_type, 16#11#),
      1618 => to_slv(opcode_type, 16#08#),
      1619 => to_slv(opcode_type, 16#06#),
      1620 => to_slv(opcode_type, 16#11#),
      1621 => to_slv(opcode_type, 16#0A#),
      1622 => to_slv(opcode_type, 16#06#),
      1623 => to_slv(opcode_type, 16#0D#),
      1624 => to_slv(opcode_type, 16#AB#),
      1625 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#08#),
      1633 => to_slv(opcode_type, 16#09#),
      1634 => to_slv(opcode_type, 16#07#),
      1635 => to_slv(opcode_type, 16#03#),
      1636 => to_slv(opcode_type, 16#0B#),
      1637 => to_slv(opcode_type, 16#08#),
      1638 => to_slv(opcode_type, 16#0F#),
      1639 => to_slv(opcode_type, 16#0D#),
      1640 => to_slv(opcode_type, 16#09#),
      1641 => to_slv(opcode_type, 16#06#),
      1642 => to_slv(opcode_type, 16#10#),
      1643 => to_slv(opcode_type, 16#0F#),
      1644 => to_slv(opcode_type, 16#01#),
      1645 => to_slv(opcode_type, 16#10#),
      1646 => to_slv(opcode_type, 16#06#),
      1647 => to_slv(opcode_type, 16#09#),
      1648 => to_slv(opcode_type, 16#06#),
      1649 => to_slv(opcode_type, 16#0C#),
      1650 => to_slv(opcode_type, 16#0C#),
      1651 => to_slv(opcode_type, 16#02#),
      1652 => to_slv(opcode_type, 16#0B#),
      1653 => to_slv(opcode_type, 16#05#),
      1654 => to_slv(opcode_type, 16#08#),
      1655 => to_slv(opcode_type, 16#0E#),
      1656 => to_slv(opcode_type, 16#0B#),
      1657 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#08#),
      1665 => to_slv(opcode_type, 16#09#),
      1666 => to_slv(opcode_type, 16#01#),
      1667 => to_slv(opcode_type, 16#01#),
      1668 => to_slv(opcode_type, 16#11#),
      1669 => to_slv(opcode_type, 16#08#),
      1670 => to_slv(opcode_type, 16#07#),
      1671 => to_slv(opcode_type, 16#0D#),
      1672 => to_slv(opcode_type, 16#0C#),
      1673 => to_slv(opcode_type, 16#06#),
      1674 => to_slv(opcode_type, 16#0B#),
      1675 => to_slv(opcode_type, 16#1C#),
      1676 => to_slv(opcode_type, 16#09#),
      1677 => to_slv(opcode_type, 16#08#),
      1678 => to_slv(opcode_type, 16#06#),
      1679 => to_slv(opcode_type, 16#0B#),
      1680 => to_slv(opcode_type, 16#0F#),
      1681 => to_slv(opcode_type, 16#05#),
      1682 => to_slv(opcode_type, 16#0B#),
      1683 => to_slv(opcode_type, 16#09#),
      1684 => to_slv(opcode_type, 16#05#),
      1685 => to_slv(opcode_type, 16#0D#),
      1686 => to_slv(opcode_type, 16#08#),
      1687 => to_slv(opcode_type, 16#0C#),
      1688 => to_slv(opcode_type, 16#0D#),
      1689 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#06#),
      1697 => to_slv(opcode_type, 16#06#),
      1698 => to_slv(opcode_type, 16#08#),
      1699 => to_slv(opcode_type, 16#03#),
      1700 => to_slv(opcode_type, 16#0A#),
      1701 => to_slv(opcode_type, 16#03#),
      1702 => to_slv(opcode_type, 16#0F#),
      1703 => to_slv(opcode_type, 16#06#),
      1704 => to_slv(opcode_type, 16#08#),
      1705 => to_slv(opcode_type, 16#11#),
      1706 => to_slv(opcode_type, 16#0C#),
      1707 => to_slv(opcode_type, 16#09#),
      1708 => to_slv(opcode_type, 16#0C#),
      1709 => to_slv(opcode_type, 16#11#),
      1710 => to_slv(opcode_type, 16#07#),
      1711 => to_slv(opcode_type, 16#01#),
      1712 => to_slv(opcode_type, 16#05#),
      1713 => to_slv(opcode_type, 16#0F#),
      1714 => to_slv(opcode_type, 16#06#),
      1715 => to_slv(opcode_type, 16#06#),
      1716 => to_slv(opcode_type, 16#0B#),
      1717 => to_slv(opcode_type, 16#0B#),
      1718 => to_slv(opcode_type, 16#06#),
      1719 => to_slv(opcode_type, 16#0A#),
      1720 => to_slv(opcode_type, 16#0B#),
      1721 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#07#),
      1729 => to_slv(opcode_type, 16#08#),
      1730 => to_slv(opcode_type, 16#01#),
      1731 => to_slv(opcode_type, 16#05#),
      1732 => to_slv(opcode_type, 16#0D#),
      1733 => to_slv(opcode_type, 16#08#),
      1734 => to_slv(opcode_type, 16#02#),
      1735 => to_slv(opcode_type, 16#0B#),
      1736 => to_slv(opcode_type, 16#05#),
      1737 => to_slv(opcode_type, 16#0E#),
      1738 => to_slv(opcode_type, 16#07#),
      1739 => to_slv(opcode_type, 16#06#),
      1740 => to_slv(opcode_type, 16#07#),
      1741 => to_slv(opcode_type, 16#0D#),
      1742 => to_slv(opcode_type, 16#0D#),
      1743 => to_slv(opcode_type, 16#07#),
      1744 => to_slv(opcode_type, 16#10#),
      1745 => to_slv(opcode_type, 16#AB#),
      1746 => to_slv(opcode_type, 16#09#),
      1747 => to_slv(opcode_type, 16#06#),
      1748 => to_slv(opcode_type, 16#0E#),
      1749 => to_slv(opcode_type, 16#0C#),
      1750 => to_slv(opcode_type, 16#07#),
      1751 => to_slv(opcode_type, 16#0B#),
      1752 => to_slv(opcode_type, 16#5F#),
      1753 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#07#),
      1761 => to_slv(opcode_type, 16#09#),
      1762 => to_slv(opcode_type, 16#04#),
      1763 => to_slv(opcode_type, 16#08#),
      1764 => to_slv(opcode_type, 16#11#),
      1765 => to_slv(opcode_type, 16#0B#),
      1766 => to_slv(opcode_type, 16#02#),
      1767 => to_slv(opcode_type, 16#09#),
      1768 => to_slv(opcode_type, 16#0E#),
      1769 => to_slv(opcode_type, 16#10#),
      1770 => to_slv(opcode_type, 16#08#),
      1771 => to_slv(opcode_type, 16#09#),
      1772 => to_slv(opcode_type, 16#07#),
      1773 => to_slv(opcode_type, 16#11#),
      1774 => to_slv(opcode_type, 16#B2#),
      1775 => to_slv(opcode_type, 16#09#),
      1776 => to_slv(opcode_type, 16#0E#),
      1777 => to_slv(opcode_type, 16#0E#),
      1778 => to_slv(opcode_type, 16#09#),
      1779 => to_slv(opcode_type, 16#08#),
      1780 => to_slv(opcode_type, 16#9B#),
      1781 => to_slv(opcode_type, 16#0D#),
      1782 => to_slv(opcode_type, 16#06#),
      1783 => to_slv(opcode_type, 16#0B#),
      1784 => to_slv(opcode_type, 16#0B#),
      1785 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#07#),
      1793 => to_slv(opcode_type, 16#06#),
      1794 => to_slv(opcode_type, 16#05#),
      1795 => to_slv(opcode_type, 16#03#),
      1796 => to_slv(opcode_type, 16#88#),
      1797 => to_slv(opcode_type, 16#09#),
      1798 => to_slv(opcode_type, 16#06#),
      1799 => to_slv(opcode_type, 16#0B#),
      1800 => to_slv(opcode_type, 16#10#),
      1801 => to_slv(opcode_type, 16#05#),
      1802 => to_slv(opcode_type, 16#0F#),
      1803 => to_slv(opcode_type, 16#07#),
      1804 => to_slv(opcode_type, 16#08#),
      1805 => to_slv(opcode_type, 16#04#),
      1806 => to_slv(opcode_type, 16#0E#),
      1807 => to_slv(opcode_type, 16#07#),
      1808 => to_slv(opcode_type, 16#CD#),
      1809 => to_slv(opcode_type, 16#11#),
      1810 => to_slv(opcode_type, 16#09#),
      1811 => to_slv(opcode_type, 16#07#),
      1812 => to_slv(opcode_type, 16#0D#),
      1813 => to_slv(opcode_type, 16#0C#),
      1814 => to_slv(opcode_type, 16#08#),
      1815 => to_slv(opcode_type, 16#0C#),
      1816 => to_slv(opcode_type, 16#0D#),
      1817 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#09#),
      1825 => to_slv(opcode_type, 16#08#),
      1826 => to_slv(opcode_type, 16#02#),
      1827 => to_slv(opcode_type, 16#02#),
      1828 => to_slv(opcode_type, 16#10#),
      1829 => to_slv(opcode_type, 16#08#),
      1830 => to_slv(opcode_type, 16#02#),
      1831 => to_slv(opcode_type, 16#0B#),
      1832 => to_slv(opcode_type, 16#05#),
      1833 => to_slv(opcode_type, 16#10#),
      1834 => to_slv(opcode_type, 16#08#),
      1835 => to_slv(opcode_type, 16#07#),
      1836 => to_slv(opcode_type, 16#08#),
      1837 => to_slv(opcode_type, 16#0F#),
      1838 => to_slv(opcode_type, 16#0B#),
      1839 => to_slv(opcode_type, 16#07#),
      1840 => to_slv(opcode_type, 16#0E#),
      1841 => to_slv(opcode_type, 16#11#),
      1842 => to_slv(opcode_type, 16#09#),
      1843 => to_slv(opcode_type, 16#07#),
      1844 => to_slv(opcode_type, 16#0B#),
      1845 => to_slv(opcode_type, 16#0B#),
      1846 => to_slv(opcode_type, 16#08#),
      1847 => to_slv(opcode_type, 16#0D#),
      1848 => to_slv(opcode_type, 16#0D#),
      1849 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#09#),
      1857 => to_slv(opcode_type, 16#07#),
      1858 => to_slv(opcode_type, 16#04#),
      1859 => to_slv(opcode_type, 16#01#),
      1860 => to_slv(opcode_type, 16#0D#),
      1861 => to_slv(opcode_type, 16#09#),
      1862 => to_slv(opcode_type, 16#08#),
      1863 => to_slv(opcode_type, 16#10#),
      1864 => to_slv(opcode_type, 16#11#),
      1865 => to_slv(opcode_type, 16#02#),
      1866 => to_slv(opcode_type, 16#0A#),
      1867 => to_slv(opcode_type, 16#07#),
      1868 => to_slv(opcode_type, 16#09#),
      1869 => to_slv(opcode_type, 16#04#),
      1870 => to_slv(opcode_type, 16#0C#),
      1871 => to_slv(opcode_type, 16#09#),
      1872 => to_slv(opcode_type, 16#0C#),
      1873 => to_slv(opcode_type, 16#10#),
      1874 => to_slv(opcode_type, 16#09#),
      1875 => to_slv(opcode_type, 16#08#),
      1876 => to_slv(opcode_type, 16#0A#),
      1877 => to_slv(opcode_type, 16#B3#),
      1878 => to_slv(opcode_type, 16#06#),
      1879 => to_slv(opcode_type, 16#0E#),
      1880 => to_slv(opcode_type, 16#0B#),
      1881 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#06#),
      1890 => to_slv(opcode_type, 16#03#),
      1891 => to_slv(opcode_type, 16#03#),
      1892 => to_slv(opcode_type, 16#11#),
      1893 => to_slv(opcode_type, 16#09#),
      1894 => to_slv(opcode_type, 16#09#),
      1895 => to_slv(opcode_type, 16#11#),
      1896 => to_slv(opcode_type, 16#11#),
      1897 => to_slv(opcode_type, 16#03#),
      1898 => to_slv(opcode_type, 16#0A#),
      1899 => to_slv(opcode_type, 16#09#),
      1900 => to_slv(opcode_type, 16#06#),
      1901 => to_slv(opcode_type, 16#08#),
      1902 => to_slv(opcode_type, 16#0A#),
      1903 => to_slv(opcode_type, 16#0C#),
      1904 => to_slv(opcode_type, 16#04#),
      1905 => to_slv(opcode_type, 16#11#),
      1906 => to_slv(opcode_type, 16#09#),
      1907 => to_slv(opcode_type, 16#06#),
      1908 => to_slv(opcode_type, 16#0A#),
      1909 => to_slv(opcode_type, 16#10#),
      1910 => to_slv(opcode_type, 16#07#),
      1911 => to_slv(opcode_type, 16#10#),
      1912 => to_slv(opcode_type, 16#0D#),
      1913 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#07#),
      1921 => to_slv(opcode_type, 16#07#),
      1922 => to_slv(opcode_type, 16#08#),
      1923 => to_slv(opcode_type, 16#01#),
      1924 => to_slv(opcode_type, 16#10#),
      1925 => to_slv(opcode_type, 16#02#),
      1926 => to_slv(opcode_type, 16#0B#),
      1927 => to_slv(opcode_type, 16#06#),
      1928 => to_slv(opcode_type, 16#02#),
      1929 => to_slv(opcode_type, 16#0E#),
      1930 => to_slv(opcode_type, 16#06#),
      1931 => to_slv(opcode_type, 16#0F#),
      1932 => to_slv(opcode_type, 16#0E#),
      1933 => to_slv(opcode_type, 16#09#),
      1934 => to_slv(opcode_type, 16#09#),
      1935 => to_slv(opcode_type, 16#08#),
      1936 => to_slv(opcode_type, 16#0E#),
      1937 => to_slv(opcode_type, 16#11#),
      1938 => to_slv(opcode_type, 16#07#),
      1939 => to_slv(opcode_type, 16#7B#),
      1940 => to_slv(opcode_type, 16#0A#),
      1941 => to_slv(opcode_type, 16#06#),
      1942 => to_slv(opcode_type, 16#04#),
      1943 => to_slv(opcode_type, 16#10#),
      1944 => to_slv(opcode_type, 16#11#),
      1945 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#08#),
      1953 => to_slv(opcode_type, 16#08#),
      1954 => to_slv(opcode_type, 16#08#),
      1955 => to_slv(opcode_type, 16#07#),
      1956 => to_slv(opcode_type, 16#C7#),
      1957 => to_slv(opcode_type, 16#0A#),
      1958 => to_slv(opcode_type, 16#03#),
      1959 => to_slv(opcode_type, 16#0C#),
      1960 => to_slv(opcode_type, 16#03#),
      1961 => to_slv(opcode_type, 16#04#),
      1962 => to_slv(opcode_type, 16#0D#),
      1963 => to_slv(opcode_type, 16#07#),
      1964 => to_slv(opcode_type, 16#08#),
      1965 => to_slv(opcode_type, 16#03#),
      1966 => to_slv(opcode_type, 16#AA#),
      1967 => to_slv(opcode_type, 16#06#),
      1968 => to_slv(opcode_type, 16#0F#),
      1969 => to_slv(opcode_type, 16#1C#),
      1970 => to_slv(opcode_type, 16#06#),
      1971 => to_slv(opcode_type, 16#09#),
      1972 => to_slv(opcode_type, 16#0D#),
      1973 => to_slv(opcode_type, 16#0C#),
      1974 => to_slv(opcode_type, 16#06#),
      1975 => to_slv(opcode_type, 16#10#),
      1976 => to_slv(opcode_type, 16#10#),
      1977 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#09#),
      1985 => to_slv(opcode_type, 16#09#),
      1986 => to_slv(opcode_type, 16#01#),
      1987 => to_slv(opcode_type, 16#09#),
      1988 => to_slv(opcode_type, 16#79#),
      1989 => to_slv(opcode_type, 16#11#),
      1990 => to_slv(opcode_type, 16#06#),
      1991 => to_slv(opcode_type, 16#01#),
      1992 => to_slv(opcode_type, 16#11#),
      1993 => to_slv(opcode_type, 16#08#),
      1994 => to_slv(opcode_type, 16#0E#),
      1995 => to_slv(opcode_type, 16#0C#),
      1996 => to_slv(opcode_type, 16#08#),
      1997 => to_slv(opcode_type, 16#06#),
      1998 => to_slv(opcode_type, 16#06#),
      1999 => to_slv(opcode_type, 16#0D#),
      2000 => to_slv(opcode_type, 16#0D#),
      2001 => to_slv(opcode_type, 16#09#),
      2002 => to_slv(opcode_type, 16#0E#),
      2003 => to_slv(opcode_type, 16#0B#),
      2004 => to_slv(opcode_type, 16#06#),
      2005 => to_slv(opcode_type, 16#04#),
      2006 => to_slv(opcode_type, 16#0C#),
      2007 => to_slv(opcode_type, 16#05#),
      2008 => to_slv(opcode_type, 16#0E#),
      2009 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#08#),
      2017 => to_slv(opcode_type, 16#09#),
      2018 => to_slv(opcode_type, 16#01#),
      2019 => to_slv(opcode_type, 16#02#),
      2020 => to_slv(opcode_type, 16#0F#),
      2021 => to_slv(opcode_type, 16#07#),
      2022 => to_slv(opcode_type, 16#04#),
      2023 => to_slv(opcode_type, 16#0E#),
      2024 => to_slv(opcode_type, 16#04#),
      2025 => to_slv(opcode_type, 16#10#),
      2026 => to_slv(opcode_type, 16#06#),
      2027 => to_slv(opcode_type, 16#06#),
      2028 => to_slv(opcode_type, 16#09#),
      2029 => to_slv(opcode_type, 16#0F#),
      2030 => to_slv(opcode_type, 16#0B#),
      2031 => to_slv(opcode_type, 16#07#),
      2032 => to_slv(opcode_type, 16#0F#),
      2033 => to_slv(opcode_type, 16#0E#),
      2034 => to_slv(opcode_type, 16#08#),
      2035 => to_slv(opcode_type, 16#08#),
      2036 => to_slv(opcode_type, 16#0B#),
      2037 => to_slv(opcode_type, 16#0B#),
      2038 => to_slv(opcode_type, 16#09#),
      2039 => to_slv(opcode_type, 16#10#),
      2040 => to_slv(opcode_type, 16#11#),
      2041 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#06#),
      2049 => to_slv(opcode_type, 16#07#),
      2050 => to_slv(opcode_type, 16#04#),
      2051 => to_slv(opcode_type, 16#08#),
      2052 => to_slv(opcode_type, 16#10#),
      2053 => to_slv(opcode_type, 16#0F#),
      2054 => to_slv(opcode_type, 16#05#),
      2055 => to_slv(opcode_type, 16#09#),
      2056 => to_slv(opcode_type, 16#0F#),
      2057 => to_slv(opcode_type, 16#10#),
      2058 => to_slv(opcode_type, 16#08#),
      2059 => to_slv(opcode_type, 16#06#),
      2060 => to_slv(opcode_type, 16#08#),
      2061 => to_slv(opcode_type, 16#0D#),
      2062 => to_slv(opcode_type, 16#11#),
      2063 => to_slv(opcode_type, 16#09#),
      2064 => to_slv(opcode_type, 16#0A#),
      2065 => to_slv(opcode_type, 16#0B#),
      2066 => to_slv(opcode_type, 16#09#),
      2067 => to_slv(opcode_type, 16#09#),
      2068 => to_slv(opcode_type, 16#0F#),
      2069 => to_slv(opcode_type, 16#11#),
      2070 => to_slv(opcode_type, 16#08#),
      2071 => to_slv(opcode_type, 16#6B#),
      2072 => to_slv(opcode_type, 16#0B#),
      2073 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#06#),
      2081 => to_slv(opcode_type, 16#09#),
      2082 => to_slv(opcode_type, 16#09#),
      2083 => to_slv(opcode_type, 16#08#),
      2084 => to_slv(opcode_type, 16#10#),
      2085 => to_slv(opcode_type, 16#0E#),
      2086 => to_slv(opcode_type, 16#05#),
      2087 => to_slv(opcode_type, 16#0B#),
      2088 => to_slv(opcode_type, 16#09#),
      2089 => to_slv(opcode_type, 16#06#),
      2090 => to_slv(opcode_type, 16#0E#),
      2091 => to_slv(opcode_type, 16#0B#),
      2092 => to_slv(opcode_type, 16#06#),
      2093 => to_slv(opcode_type, 16#55#),
      2094 => to_slv(opcode_type, 16#0E#),
      2095 => to_slv(opcode_type, 16#09#),
      2096 => to_slv(opcode_type, 16#08#),
      2097 => to_slv(opcode_type, 16#03#),
      2098 => to_slv(opcode_type, 16#0F#),
      2099 => to_slv(opcode_type, 16#03#),
      2100 => to_slv(opcode_type, 16#0A#),
      2101 => to_slv(opcode_type, 16#06#),
      2102 => to_slv(opcode_type, 16#04#),
      2103 => to_slv(opcode_type, 16#11#),
      2104 => to_slv(opcode_type, 16#0B#),
      2105 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#07#),
      2113 => to_slv(opcode_type, 16#09#),
      2114 => to_slv(opcode_type, 16#08#),
      2115 => to_slv(opcode_type, 16#01#),
      2116 => to_slv(opcode_type, 16#0A#),
      2117 => to_slv(opcode_type, 16#03#),
      2118 => to_slv(opcode_type, 16#0B#),
      2119 => to_slv(opcode_type, 16#09#),
      2120 => to_slv(opcode_type, 16#05#),
      2121 => to_slv(opcode_type, 16#0F#),
      2122 => to_slv(opcode_type, 16#07#),
      2123 => to_slv(opcode_type, 16#10#),
      2124 => to_slv(opcode_type, 16#11#),
      2125 => to_slv(opcode_type, 16#06#),
      2126 => to_slv(opcode_type, 16#05#),
      2127 => to_slv(opcode_type, 16#07#),
      2128 => to_slv(opcode_type, 16#0B#),
      2129 => to_slv(opcode_type, 16#11#),
      2130 => to_slv(opcode_type, 16#06#),
      2131 => to_slv(opcode_type, 16#06#),
      2132 => to_slv(opcode_type, 16#0E#),
      2133 => to_slv(opcode_type, 16#11#),
      2134 => to_slv(opcode_type, 16#07#),
      2135 => to_slv(opcode_type, 16#98#),
      2136 => to_slv(opcode_type, 16#0F#),
      2137 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#08#),
      2146 => to_slv(opcode_type, 16#03#),
      2147 => to_slv(opcode_type, 16#08#),
      2148 => to_slv(opcode_type, 16#0F#),
      2149 => to_slv(opcode_type, 16#0C#),
      2150 => to_slv(opcode_type, 16#09#),
      2151 => to_slv(opcode_type, 16#07#),
      2152 => to_slv(opcode_type, 16#0B#),
      2153 => to_slv(opcode_type, 16#0C#),
      2154 => to_slv(opcode_type, 16#07#),
      2155 => to_slv(opcode_type, 16#0D#),
      2156 => to_slv(opcode_type, 16#10#),
      2157 => to_slv(opcode_type, 16#07#),
      2158 => to_slv(opcode_type, 16#02#),
      2159 => to_slv(opcode_type, 16#06#),
      2160 => to_slv(opcode_type, 16#0E#),
      2161 => to_slv(opcode_type, 16#0B#),
      2162 => to_slv(opcode_type, 16#06#),
      2163 => to_slv(opcode_type, 16#08#),
      2164 => to_slv(opcode_type, 16#0D#),
      2165 => to_slv(opcode_type, 16#0A#),
      2166 => to_slv(opcode_type, 16#09#),
      2167 => to_slv(opcode_type, 16#11#),
      2168 => to_slv(opcode_type, 16#0D#),
      2169 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#09#),
      2177 => to_slv(opcode_type, 16#09#),
      2178 => to_slv(opcode_type, 16#06#),
      2179 => to_slv(opcode_type, 16#07#),
      2180 => to_slv(opcode_type, 16#0F#),
      2181 => to_slv(opcode_type, 16#0B#),
      2182 => to_slv(opcode_type, 16#02#),
      2183 => to_slv(opcode_type, 16#0C#),
      2184 => to_slv(opcode_type, 16#08#),
      2185 => to_slv(opcode_type, 16#05#),
      2186 => to_slv(opcode_type, 16#0D#),
      2187 => to_slv(opcode_type, 16#06#),
      2188 => to_slv(opcode_type, 16#0B#),
      2189 => to_slv(opcode_type, 16#0A#),
      2190 => to_slv(opcode_type, 16#06#),
      2191 => to_slv(opcode_type, 16#05#),
      2192 => to_slv(opcode_type, 16#07#),
      2193 => to_slv(opcode_type, 16#10#),
      2194 => to_slv(opcode_type, 16#0E#),
      2195 => to_slv(opcode_type, 16#09#),
      2196 => to_slv(opcode_type, 16#09#),
      2197 => to_slv(opcode_type, 16#0B#),
      2198 => to_slv(opcode_type, 16#0F#),
      2199 => to_slv(opcode_type, 16#03#),
      2200 => to_slv(opcode_type, 16#0F#),
      2201 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#07#),
      2209 => to_slv(opcode_type, 16#09#),
      2210 => to_slv(opcode_type, 16#03#),
      2211 => to_slv(opcode_type, 16#07#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#0F#),
      2214 => to_slv(opcode_type, 16#02#),
      2215 => to_slv(opcode_type, 16#08#),
      2216 => to_slv(opcode_type, 16#0C#),
      2217 => to_slv(opcode_type, 16#0F#),
      2218 => to_slv(opcode_type, 16#06#),
      2219 => to_slv(opcode_type, 16#08#),
      2220 => to_slv(opcode_type, 16#08#),
      2221 => to_slv(opcode_type, 16#0E#),
      2222 => to_slv(opcode_type, 16#0A#),
      2223 => to_slv(opcode_type, 16#08#),
      2224 => to_slv(opcode_type, 16#0B#),
      2225 => to_slv(opcode_type, 16#0F#),
      2226 => to_slv(opcode_type, 16#08#),
      2227 => to_slv(opcode_type, 16#07#),
      2228 => to_slv(opcode_type, 16#0A#),
      2229 => to_slv(opcode_type, 16#10#),
      2230 => to_slv(opcode_type, 16#06#),
      2231 => to_slv(opcode_type, 16#11#),
      2232 => to_slv(opcode_type, 16#10#),
      2233 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#06#),
      2242 => to_slv(opcode_type, 16#03#),
      2243 => to_slv(opcode_type, 16#08#),
      2244 => to_slv(opcode_type, 16#10#),
      2245 => to_slv(opcode_type, 16#10#),
      2246 => to_slv(opcode_type, 16#02#),
      2247 => to_slv(opcode_type, 16#06#),
      2248 => to_slv(opcode_type, 16#0E#),
      2249 => to_slv(opcode_type, 16#0F#),
      2250 => to_slv(opcode_type, 16#09#),
      2251 => to_slv(opcode_type, 16#08#),
      2252 => to_slv(opcode_type, 16#07#),
      2253 => to_slv(opcode_type, 16#0E#),
      2254 => to_slv(opcode_type, 16#0B#),
      2255 => to_slv(opcode_type, 16#06#),
      2256 => to_slv(opcode_type, 16#11#),
      2257 => to_slv(opcode_type, 16#0C#),
      2258 => to_slv(opcode_type, 16#09#),
      2259 => to_slv(opcode_type, 16#09#),
      2260 => to_slv(opcode_type, 16#0C#),
      2261 => to_slv(opcode_type, 16#0B#),
      2262 => to_slv(opcode_type, 16#07#),
      2263 => to_slv(opcode_type, 16#11#),
      2264 => to_slv(opcode_type, 16#0F#),
      2265 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#06#),
      2273 => to_slv(opcode_type, 16#06#),
      2274 => to_slv(opcode_type, 16#09#),
      2275 => to_slv(opcode_type, 16#05#),
      2276 => to_slv(opcode_type, 16#11#),
      2277 => to_slv(opcode_type, 16#07#),
      2278 => to_slv(opcode_type, 16#0E#),
      2279 => to_slv(opcode_type, 16#11#),
      2280 => to_slv(opcode_type, 16#03#),
      2281 => to_slv(opcode_type, 16#02#),
      2282 => to_slv(opcode_type, 16#0D#),
      2283 => to_slv(opcode_type, 16#08#),
      2284 => to_slv(opcode_type, 16#09#),
      2285 => to_slv(opcode_type, 16#04#),
      2286 => to_slv(opcode_type, 16#0A#),
      2287 => to_slv(opcode_type, 16#08#),
      2288 => to_slv(opcode_type, 16#0C#),
      2289 => to_slv(opcode_type, 16#0D#),
      2290 => to_slv(opcode_type, 16#08#),
      2291 => to_slv(opcode_type, 16#08#),
      2292 => to_slv(opcode_type, 16#99#),
      2293 => to_slv(opcode_type, 16#0A#),
      2294 => to_slv(opcode_type, 16#08#),
      2295 => to_slv(opcode_type, 16#0D#),
      2296 => to_slv(opcode_type, 16#0A#),
      2297 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#09#),
      2305 => to_slv(opcode_type, 16#07#),
      2306 => to_slv(opcode_type, 16#05#),
      2307 => to_slv(opcode_type, 16#06#),
      2308 => to_slv(opcode_type, 16#0E#),
      2309 => to_slv(opcode_type, 16#11#),
      2310 => to_slv(opcode_type, 16#07#),
      2311 => to_slv(opcode_type, 16#07#),
      2312 => to_slv(opcode_type, 16#0A#),
      2313 => to_slv(opcode_type, 16#10#),
      2314 => to_slv(opcode_type, 16#03#),
      2315 => to_slv(opcode_type, 16#0F#),
      2316 => to_slv(opcode_type, 16#08#),
      2317 => to_slv(opcode_type, 16#09#),
      2318 => to_slv(opcode_type, 16#05#),
      2319 => to_slv(opcode_type, 16#0B#),
      2320 => to_slv(opcode_type, 16#01#),
      2321 => to_slv(opcode_type, 16#0F#),
      2322 => to_slv(opcode_type, 16#06#),
      2323 => to_slv(opcode_type, 16#07#),
      2324 => to_slv(opcode_type, 16#0B#),
      2325 => to_slv(opcode_type, 16#0B#),
      2326 => to_slv(opcode_type, 16#07#),
      2327 => to_slv(opcode_type, 16#0C#),
      2328 => to_slv(opcode_type, 16#0D#),
      2329 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#09#),
      2337 => to_slv(opcode_type, 16#06#),
      2338 => to_slv(opcode_type, 16#01#),
      2339 => to_slv(opcode_type, 16#09#),
      2340 => to_slv(opcode_type, 16#0B#),
      2341 => to_slv(opcode_type, 16#10#),
      2342 => to_slv(opcode_type, 16#09#),
      2343 => to_slv(opcode_type, 16#02#),
      2344 => to_slv(opcode_type, 16#0D#),
      2345 => to_slv(opcode_type, 16#05#),
      2346 => to_slv(opcode_type, 16#11#),
      2347 => to_slv(opcode_type, 16#09#),
      2348 => to_slv(opcode_type, 16#06#),
      2349 => to_slv(opcode_type, 16#02#),
      2350 => to_slv(opcode_type, 16#0A#),
      2351 => to_slv(opcode_type, 16#08#),
      2352 => to_slv(opcode_type, 16#0E#),
      2353 => to_slv(opcode_type, 16#0F#),
      2354 => to_slv(opcode_type, 16#08#),
      2355 => to_slv(opcode_type, 16#09#),
      2356 => to_slv(opcode_type, 16#10#),
      2357 => to_slv(opcode_type, 16#11#),
      2358 => to_slv(opcode_type, 16#08#),
      2359 => to_slv(opcode_type, 16#11#),
      2360 => to_slv(opcode_type, 16#0D#),
      2361 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#09#),
      2369 => to_slv(opcode_type, 16#06#),
      2370 => to_slv(opcode_type, 16#01#),
      2371 => to_slv(opcode_type, 16#05#),
      2372 => to_slv(opcode_type, 16#0C#),
      2373 => to_slv(opcode_type, 16#08#),
      2374 => to_slv(opcode_type, 16#06#),
      2375 => to_slv(opcode_type, 16#10#),
      2376 => to_slv(opcode_type, 16#0C#),
      2377 => to_slv(opcode_type, 16#06#),
      2378 => to_slv(opcode_type, 16#10#),
      2379 => to_slv(opcode_type, 16#0B#),
      2380 => to_slv(opcode_type, 16#09#),
      2381 => to_slv(opcode_type, 16#09#),
      2382 => to_slv(opcode_type, 16#01#),
      2383 => to_slv(opcode_type, 16#10#),
      2384 => to_slv(opcode_type, 16#03#),
      2385 => to_slv(opcode_type, 16#0E#),
      2386 => to_slv(opcode_type, 16#06#),
      2387 => to_slv(opcode_type, 16#09#),
      2388 => to_slv(opcode_type, 16#10#),
      2389 => to_slv(opcode_type, 16#0E#),
      2390 => to_slv(opcode_type, 16#06#),
      2391 => to_slv(opcode_type, 16#0F#),
      2392 => to_slv(opcode_type, 16#0B#),
      2393 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#07#),
      2402 => to_slv(opcode_type, 16#08#),
      2403 => to_slv(opcode_type, 16#02#),
      2404 => to_slv(opcode_type, 16#0D#),
      2405 => to_slv(opcode_type, 16#06#),
      2406 => to_slv(opcode_type, 16#0B#),
      2407 => to_slv(opcode_type, 16#11#),
      2408 => to_slv(opcode_type, 16#09#),
      2409 => to_slv(opcode_type, 16#02#),
      2410 => to_slv(opcode_type, 16#2E#),
      2411 => to_slv(opcode_type, 16#04#),
      2412 => to_slv(opcode_type, 16#10#),
      2413 => to_slv(opcode_type, 16#08#),
      2414 => to_slv(opcode_type, 16#08#),
      2415 => to_slv(opcode_type, 16#02#),
      2416 => to_slv(opcode_type, 16#11#),
      2417 => to_slv(opcode_type, 16#06#),
      2418 => to_slv(opcode_type, 16#10#),
      2419 => to_slv(opcode_type, 16#10#),
      2420 => to_slv(opcode_type, 16#07#),
      2421 => to_slv(opcode_type, 16#04#),
      2422 => to_slv(opcode_type, 16#BD#),
      2423 => to_slv(opcode_type, 16#05#),
      2424 => to_slv(opcode_type, 16#11#),
      2425 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#09#),
      2433 => to_slv(opcode_type, 16#06#),
      2434 => to_slv(opcode_type, 16#01#),
      2435 => to_slv(opcode_type, 16#03#),
      2436 => to_slv(opcode_type, 16#0F#),
      2437 => to_slv(opcode_type, 16#06#),
      2438 => to_slv(opcode_type, 16#03#),
      2439 => to_slv(opcode_type, 16#68#),
      2440 => to_slv(opcode_type, 16#01#),
      2441 => to_slv(opcode_type, 16#0B#),
      2442 => to_slv(opcode_type, 16#06#),
      2443 => to_slv(opcode_type, 16#06#),
      2444 => to_slv(opcode_type, 16#08#),
      2445 => to_slv(opcode_type, 16#0C#),
      2446 => to_slv(opcode_type, 16#CD#),
      2447 => to_slv(opcode_type, 16#07#),
      2448 => to_slv(opcode_type, 16#6B#),
      2449 => to_slv(opcode_type, 16#11#),
      2450 => to_slv(opcode_type, 16#06#),
      2451 => to_slv(opcode_type, 16#09#),
      2452 => to_slv(opcode_type, 16#D9#),
      2453 => to_slv(opcode_type, 16#25#),
      2454 => to_slv(opcode_type, 16#06#),
      2455 => to_slv(opcode_type, 16#0A#),
      2456 => to_slv(opcode_type, 16#0A#),
      2457 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#07#),
      2465 => to_slv(opcode_type, 16#07#),
      2466 => to_slv(opcode_type, 16#02#),
      2467 => to_slv(opcode_type, 16#08#),
      2468 => to_slv(opcode_type, 16#0E#),
      2469 => to_slv(opcode_type, 16#11#),
      2470 => to_slv(opcode_type, 16#04#),
      2471 => to_slv(opcode_type, 16#06#),
      2472 => to_slv(opcode_type, 16#0C#),
      2473 => to_slv(opcode_type, 16#B2#),
      2474 => to_slv(opcode_type, 16#06#),
      2475 => to_slv(opcode_type, 16#07#),
      2476 => to_slv(opcode_type, 16#06#),
      2477 => to_slv(opcode_type, 16#0E#),
      2478 => to_slv(opcode_type, 16#1C#),
      2479 => to_slv(opcode_type, 16#06#),
      2480 => to_slv(opcode_type, 16#CC#),
      2481 => to_slv(opcode_type, 16#A5#),
      2482 => to_slv(opcode_type, 16#08#),
      2483 => to_slv(opcode_type, 16#06#),
      2484 => to_slv(opcode_type, 16#0D#),
      2485 => to_slv(opcode_type, 16#0A#),
      2486 => to_slv(opcode_type, 16#09#),
      2487 => to_slv(opcode_type, 16#0F#),
      2488 => to_slv(opcode_type, 16#C1#),
      2489 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#07#),
      2497 => to_slv(opcode_type, 16#08#),
      2498 => to_slv(opcode_type, 16#09#),
      2499 => to_slv(opcode_type, 16#06#),
      2500 => to_slv(opcode_type, 16#0A#),
      2501 => to_slv(opcode_type, 16#0A#),
      2502 => to_slv(opcode_type, 16#05#),
      2503 => to_slv(opcode_type, 16#10#),
      2504 => to_slv(opcode_type, 16#07#),
      2505 => to_slv(opcode_type, 16#02#),
      2506 => to_slv(opcode_type, 16#27#),
      2507 => to_slv(opcode_type, 16#03#),
      2508 => to_slv(opcode_type, 16#0B#),
      2509 => to_slv(opcode_type, 16#08#),
      2510 => to_slv(opcode_type, 16#04#),
      2511 => to_slv(opcode_type, 16#06#),
      2512 => to_slv(opcode_type, 16#10#),
      2513 => to_slv(opcode_type, 16#0B#),
      2514 => to_slv(opcode_type, 16#07#),
      2515 => to_slv(opcode_type, 16#08#),
      2516 => to_slv(opcode_type, 16#0B#),
      2517 => to_slv(opcode_type, 16#0A#),
      2518 => to_slv(opcode_type, 16#08#),
      2519 => to_slv(opcode_type, 16#E5#),
      2520 => to_slv(opcode_type, 16#0A#),
      2521 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#07#),
      2530 => to_slv(opcode_type, 16#08#),
      2531 => to_slv(opcode_type, 16#04#),
      2532 => to_slv(opcode_type, 16#CA#),
      2533 => to_slv(opcode_type, 16#03#),
      2534 => to_slv(opcode_type, 16#11#),
      2535 => to_slv(opcode_type, 16#01#),
      2536 => to_slv(opcode_type, 16#07#),
      2537 => to_slv(opcode_type, 16#11#),
      2538 => to_slv(opcode_type, 16#0D#),
      2539 => to_slv(opcode_type, 16#08#),
      2540 => to_slv(opcode_type, 16#08#),
      2541 => to_slv(opcode_type, 16#03#),
      2542 => to_slv(opcode_type, 16#0F#),
      2543 => to_slv(opcode_type, 16#09#),
      2544 => to_slv(opcode_type, 16#0A#),
      2545 => to_slv(opcode_type, 16#0A#),
      2546 => to_slv(opcode_type, 16#07#),
      2547 => to_slv(opcode_type, 16#07#),
      2548 => to_slv(opcode_type, 16#0B#),
      2549 => to_slv(opcode_type, 16#10#),
      2550 => to_slv(opcode_type, 16#07#),
      2551 => to_slv(opcode_type, 16#D0#),
      2552 => to_slv(opcode_type, 16#0B#),
      2553 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#07#),
      2561 => to_slv(opcode_type, 16#07#),
      2562 => to_slv(opcode_type, 16#07#),
      2563 => to_slv(opcode_type, 16#05#),
      2564 => to_slv(opcode_type, 16#EB#),
      2565 => to_slv(opcode_type, 16#07#),
      2566 => to_slv(opcode_type, 16#0C#),
      2567 => to_slv(opcode_type, 16#0D#),
      2568 => to_slv(opcode_type, 16#01#),
      2569 => to_slv(opcode_type, 16#04#),
      2570 => to_slv(opcode_type, 16#10#),
      2571 => to_slv(opcode_type, 16#08#),
      2572 => to_slv(opcode_type, 16#07#),
      2573 => to_slv(opcode_type, 16#09#),
      2574 => to_slv(opcode_type, 16#0A#),
      2575 => to_slv(opcode_type, 16#0F#),
      2576 => to_slv(opcode_type, 16#09#),
      2577 => to_slv(opcode_type, 16#10#),
      2578 => to_slv(opcode_type, 16#0A#),
      2579 => to_slv(opcode_type, 16#06#),
      2580 => to_slv(opcode_type, 16#02#),
      2581 => to_slv(opcode_type, 16#11#),
      2582 => to_slv(opcode_type, 16#07#),
      2583 => to_slv(opcode_type, 16#0D#),
      2584 => to_slv(opcode_type, 16#0B#),
      2585 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#06#),
      2593 => to_slv(opcode_type, 16#07#),
      2594 => to_slv(opcode_type, 16#04#),
      2595 => to_slv(opcode_type, 16#01#),
      2596 => to_slv(opcode_type, 16#0A#),
      2597 => to_slv(opcode_type, 16#07#),
      2598 => to_slv(opcode_type, 16#01#),
      2599 => to_slv(opcode_type, 16#0D#),
      2600 => to_slv(opcode_type, 16#07#),
      2601 => to_slv(opcode_type, 16#0F#),
      2602 => to_slv(opcode_type, 16#0E#),
      2603 => to_slv(opcode_type, 16#09#),
      2604 => to_slv(opcode_type, 16#09#),
      2605 => to_slv(opcode_type, 16#08#),
      2606 => to_slv(opcode_type, 16#0F#),
      2607 => to_slv(opcode_type, 16#0E#),
      2608 => to_slv(opcode_type, 16#03#),
      2609 => to_slv(opcode_type, 16#11#),
      2610 => to_slv(opcode_type, 16#09#),
      2611 => to_slv(opcode_type, 16#07#),
      2612 => to_slv(opcode_type, 16#0A#),
      2613 => to_slv(opcode_type, 16#87#),
      2614 => to_slv(opcode_type, 16#09#),
      2615 => to_slv(opcode_type, 16#0D#),
      2616 => to_slv(opcode_type, 16#0C#),
      2617 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#07#),
      2625 => to_slv(opcode_type, 16#09#),
      2626 => to_slv(opcode_type, 16#06#),
      2627 => to_slv(opcode_type, 16#01#),
      2628 => to_slv(opcode_type, 16#0E#),
      2629 => to_slv(opcode_type, 16#01#),
      2630 => to_slv(opcode_type, 16#0E#),
      2631 => to_slv(opcode_type, 16#07#),
      2632 => to_slv(opcode_type, 16#06#),
      2633 => to_slv(opcode_type, 16#0B#),
      2634 => to_slv(opcode_type, 16#11#),
      2635 => to_slv(opcode_type, 16#09#),
      2636 => to_slv(opcode_type, 16#0D#),
      2637 => to_slv(opcode_type, 16#0A#),
      2638 => to_slv(opcode_type, 16#07#),
      2639 => to_slv(opcode_type, 16#07#),
      2640 => to_slv(opcode_type, 16#08#),
      2641 => to_slv(opcode_type, 16#53#),
      2642 => to_slv(opcode_type, 16#10#),
      2643 => to_slv(opcode_type, 16#04#),
      2644 => to_slv(opcode_type, 16#0E#),
      2645 => to_slv(opcode_type, 16#03#),
      2646 => to_slv(opcode_type, 16#08#),
      2647 => to_slv(opcode_type, 16#0C#),
      2648 => to_slv(opcode_type, 16#0C#),
      2649 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#09#),
      2657 => to_slv(opcode_type, 16#07#),
      2658 => to_slv(opcode_type, 16#04#),
      2659 => to_slv(opcode_type, 16#01#),
      2660 => to_slv(opcode_type, 16#0E#),
      2661 => to_slv(opcode_type, 16#09#),
      2662 => to_slv(opcode_type, 16#02#),
      2663 => to_slv(opcode_type, 16#0B#),
      2664 => to_slv(opcode_type, 16#02#),
      2665 => to_slv(opcode_type, 16#11#),
      2666 => to_slv(opcode_type, 16#08#),
      2667 => to_slv(opcode_type, 16#07#),
      2668 => to_slv(opcode_type, 16#09#),
      2669 => to_slv(opcode_type, 16#0E#),
      2670 => to_slv(opcode_type, 16#0E#),
      2671 => to_slv(opcode_type, 16#09#),
      2672 => to_slv(opcode_type, 16#47#),
      2673 => to_slv(opcode_type, 16#0F#),
      2674 => to_slv(opcode_type, 16#06#),
      2675 => to_slv(opcode_type, 16#06#),
      2676 => to_slv(opcode_type, 16#0A#),
      2677 => to_slv(opcode_type, 16#0C#),
      2678 => to_slv(opcode_type, 16#06#),
      2679 => to_slv(opcode_type, 16#10#),
      2680 => to_slv(opcode_type, 16#0B#),
      2681 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#06#),
      2689 => to_slv(opcode_type, 16#09#),
      2690 => to_slv(opcode_type, 16#01#),
      2691 => to_slv(opcode_type, 16#03#),
      2692 => to_slv(opcode_type, 16#8E#),
      2693 => to_slv(opcode_type, 16#06#),
      2694 => to_slv(opcode_type, 16#09#),
      2695 => to_slv(opcode_type, 16#10#),
      2696 => to_slv(opcode_type, 16#18#),
      2697 => to_slv(opcode_type, 16#03#),
      2698 => to_slv(opcode_type, 16#0B#),
      2699 => to_slv(opcode_type, 16#08#),
      2700 => to_slv(opcode_type, 16#09#),
      2701 => to_slv(opcode_type, 16#07#),
      2702 => to_slv(opcode_type, 16#0B#),
      2703 => to_slv(opcode_type, 16#0C#),
      2704 => to_slv(opcode_type, 16#06#),
      2705 => to_slv(opcode_type, 16#0F#),
      2706 => to_slv(opcode_type, 16#10#),
      2707 => to_slv(opcode_type, 16#07#),
      2708 => to_slv(opcode_type, 16#09#),
      2709 => to_slv(opcode_type, 16#0A#),
      2710 => to_slv(opcode_type, 16#0B#),
      2711 => to_slv(opcode_type, 16#01#),
      2712 => to_slv(opcode_type, 16#0A#),
      2713 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#07#),
      2721 => to_slv(opcode_type, 16#06#),
      2722 => to_slv(opcode_type, 16#08#),
      2723 => to_slv(opcode_type, 16#04#),
      2724 => to_slv(opcode_type, 16#0D#),
      2725 => to_slv(opcode_type, 16#08#),
      2726 => to_slv(opcode_type, 16#0C#),
      2727 => to_slv(opcode_type, 16#0F#),
      2728 => to_slv(opcode_type, 16#08#),
      2729 => to_slv(opcode_type, 16#01#),
      2730 => to_slv(opcode_type, 16#0F#),
      2731 => to_slv(opcode_type, 16#05#),
      2732 => to_slv(opcode_type, 16#0D#),
      2733 => to_slv(opcode_type, 16#08#),
      2734 => to_slv(opcode_type, 16#01#),
      2735 => to_slv(opcode_type, 16#06#),
      2736 => to_slv(opcode_type, 16#0B#),
      2737 => to_slv(opcode_type, 16#10#),
      2738 => to_slv(opcode_type, 16#08#),
      2739 => to_slv(opcode_type, 16#08#),
      2740 => to_slv(opcode_type, 16#0E#),
      2741 => to_slv(opcode_type, 16#24#),
      2742 => to_slv(opcode_type, 16#06#),
      2743 => to_slv(opcode_type, 16#10#),
      2744 => to_slv(opcode_type, 16#0D#),
      2745 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#07#),
      2753 => to_slv(opcode_type, 16#09#),
      2754 => to_slv(opcode_type, 16#08#),
      2755 => to_slv(opcode_type, 16#06#),
      2756 => to_slv(opcode_type, 16#11#),
      2757 => to_slv(opcode_type, 16#A6#),
      2758 => to_slv(opcode_type, 16#09#),
      2759 => to_slv(opcode_type, 16#0A#),
      2760 => to_slv(opcode_type, 16#10#),
      2761 => to_slv(opcode_type, 16#03#),
      2762 => to_slv(opcode_type, 16#01#),
      2763 => to_slv(opcode_type, 16#0F#),
      2764 => to_slv(opcode_type, 16#06#),
      2765 => to_slv(opcode_type, 16#07#),
      2766 => to_slv(opcode_type, 16#08#),
      2767 => to_slv(opcode_type, 16#10#),
      2768 => to_slv(opcode_type, 16#0E#),
      2769 => to_slv(opcode_type, 16#04#),
      2770 => to_slv(opcode_type, 16#0C#),
      2771 => to_slv(opcode_type, 16#07#),
      2772 => to_slv(opcode_type, 16#03#),
      2773 => to_slv(opcode_type, 16#0F#),
      2774 => to_slv(opcode_type, 16#09#),
      2775 => to_slv(opcode_type, 16#0D#),
      2776 => to_slv(opcode_type, 16#0D#),
      2777 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#06#),
      2785 => to_slv(opcode_type, 16#09#),
      2786 => to_slv(opcode_type, 16#04#),
      2787 => to_slv(opcode_type, 16#08#),
      2788 => to_slv(opcode_type, 16#0D#),
      2789 => to_slv(opcode_type, 16#0C#),
      2790 => to_slv(opcode_type, 16#04#),
      2791 => to_slv(opcode_type, 16#07#),
      2792 => to_slv(opcode_type, 16#13#),
      2793 => to_slv(opcode_type, 16#0C#),
      2794 => to_slv(opcode_type, 16#06#),
      2795 => to_slv(opcode_type, 16#06#),
      2796 => to_slv(opcode_type, 16#06#),
      2797 => to_slv(opcode_type, 16#0D#),
      2798 => to_slv(opcode_type, 16#0E#),
      2799 => to_slv(opcode_type, 16#09#),
      2800 => to_slv(opcode_type, 16#10#),
      2801 => to_slv(opcode_type, 16#0E#),
      2802 => to_slv(opcode_type, 16#08#),
      2803 => to_slv(opcode_type, 16#08#),
      2804 => to_slv(opcode_type, 16#0E#),
      2805 => to_slv(opcode_type, 16#F2#),
      2806 => to_slv(opcode_type, 16#07#),
      2807 => to_slv(opcode_type, 16#0C#),
      2808 => to_slv(opcode_type, 16#0B#),
      2809 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#07#),
      2817 => to_slv(opcode_type, 16#08#),
      2818 => to_slv(opcode_type, 16#08#),
      2819 => to_slv(opcode_type, 16#07#),
      2820 => to_slv(opcode_type, 16#0E#),
      2821 => to_slv(opcode_type, 16#0C#),
      2822 => to_slv(opcode_type, 16#06#),
      2823 => to_slv(opcode_type, 16#EC#),
      2824 => to_slv(opcode_type, 16#0A#),
      2825 => to_slv(opcode_type, 16#04#),
      2826 => to_slv(opcode_type, 16#01#),
      2827 => to_slv(opcode_type, 16#60#),
      2828 => to_slv(opcode_type, 16#08#),
      2829 => to_slv(opcode_type, 16#09#),
      2830 => to_slv(opcode_type, 16#09#),
      2831 => to_slv(opcode_type, 16#0F#),
      2832 => to_slv(opcode_type, 16#0F#),
      2833 => to_slv(opcode_type, 16#01#),
      2834 => to_slv(opcode_type, 16#80#),
      2835 => to_slv(opcode_type, 16#06#),
      2836 => to_slv(opcode_type, 16#07#),
      2837 => to_slv(opcode_type, 16#10#),
      2838 => to_slv(opcode_type, 16#11#),
      2839 => to_slv(opcode_type, 16#05#),
      2840 => to_slv(opcode_type, 16#0E#),
      2841 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#08#),
      2849 => to_slv(opcode_type, 16#07#),
      2850 => to_slv(opcode_type, 16#02#),
      2851 => to_slv(opcode_type, 16#09#),
      2852 => to_slv(opcode_type, 16#CA#),
      2853 => to_slv(opcode_type, 16#0D#),
      2854 => to_slv(opcode_type, 16#08#),
      2855 => to_slv(opcode_type, 16#01#),
      2856 => to_slv(opcode_type, 16#10#),
      2857 => to_slv(opcode_type, 16#02#),
      2858 => to_slv(opcode_type, 16#0D#),
      2859 => to_slv(opcode_type, 16#06#),
      2860 => to_slv(opcode_type, 16#09#),
      2861 => to_slv(opcode_type, 16#01#),
      2862 => to_slv(opcode_type, 16#0F#),
      2863 => to_slv(opcode_type, 16#07#),
      2864 => to_slv(opcode_type, 16#0F#),
      2865 => to_slv(opcode_type, 16#0B#),
      2866 => to_slv(opcode_type, 16#06#),
      2867 => to_slv(opcode_type, 16#06#),
      2868 => to_slv(opcode_type, 16#10#),
      2869 => to_slv(opcode_type, 16#0F#),
      2870 => to_slv(opcode_type, 16#08#),
      2871 => to_slv(opcode_type, 16#71#),
      2872 => to_slv(opcode_type, 16#0D#),
      2873 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#08#),
      2881 => to_slv(opcode_type, 16#06#),
      2882 => to_slv(opcode_type, 16#07#),
      2883 => to_slv(opcode_type, 16#07#),
      2884 => to_slv(opcode_type, 16#0F#),
      2885 => to_slv(opcode_type, 16#0D#),
      2886 => to_slv(opcode_type, 16#02#),
      2887 => to_slv(opcode_type, 16#20#),
      2888 => to_slv(opcode_type, 16#04#),
      2889 => to_slv(opcode_type, 16#01#),
      2890 => to_slv(opcode_type, 16#0B#),
      2891 => to_slv(opcode_type, 16#08#),
      2892 => to_slv(opcode_type, 16#08#),
      2893 => to_slv(opcode_type, 16#05#),
      2894 => to_slv(opcode_type, 16#0C#),
      2895 => to_slv(opcode_type, 16#07#),
      2896 => to_slv(opcode_type, 16#11#),
      2897 => to_slv(opcode_type, 16#11#),
      2898 => to_slv(opcode_type, 16#08#),
      2899 => to_slv(opcode_type, 16#07#),
      2900 => to_slv(opcode_type, 16#0C#),
      2901 => to_slv(opcode_type, 16#0D#),
      2902 => to_slv(opcode_type, 16#09#),
      2903 => to_slv(opcode_type, 16#0D#),
      2904 => to_slv(opcode_type, 16#0F#),
      2905 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#08#),
      2913 => to_slv(opcode_type, 16#09#),
      2914 => to_slv(opcode_type, 16#06#),
      2915 => to_slv(opcode_type, 16#06#),
      2916 => to_slv(opcode_type, 16#0C#),
      2917 => to_slv(opcode_type, 16#0E#),
      2918 => to_slv(opcode_type, 16#01#),
      2919 => to_slv(opcode_type, 16#0A#),
      2920 => to_slv(opcode_type, 16#08#),
      2921 => to_slv(opcode_type, 16#08#),
      2922 => to_slv(opcode_type, 16#10#),
      2923 => to_slv(opcode_type, 16#0E#),
      2924 => to_slv(opcode_type, 16#02#),
      2925 => to_slv(opcode_type, 16#0A#),
      2926 => to_slv(opcode_type, 16#08#),
      2927 => to_slv(opcode_type, 16#01#),
      2928 => to_slv(opcode_type, 16#05#),
      2929 => to_slv(opcode_type, 16#6A#),
      2930 => to_slv(opcode_type, 16#08#),
      2931 => to_slv(opcode_type, 16#06#),
      2932 => to_slv(opcode_type, 16#0F#),
      2933 => to_slv(opcode_type, 16#0B#),
      2934 => to_slv(opcode_type, 16#07#),
      2935 => to_slv(opcode_type, 16#10#),
      2936 => to_slv(opcode_type, 16#0D#),
      2937 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#07#),
      2945 => to_slv(opcode_type, 16#06#),
      2946 => to_slv(opcode_type, 16#04#),
      2947 => to_slv(opcode_type, 16#03#),
      2948 => to_slv(opcode_type, 16#0A#),
      2949 => to_slv(opcode_type, 16#08#),
      2950 => to_slv(opcode_type, 16#02#),
      2951 => to_slv(opcode_type, 16#0E#),
      2952 => to_slv(opcode_type, 16#07#),
      2953 => to_slv(opcode_type, 16#A8#),
      2954 => to_slv(opcode_type, 16#0B#),
      2955 => to_slv(opcode_type, 16#06#),
      2956 => to_slv(opcode_type, 16#07#),
      2957 => to_slv(opcode_type, 16#09#),
      2958 => to_slv(opcode_type, 16#0A#),
      2959 => to_slv(opcode_type, 16#0F#),
      2960 => to_slv(opcode_type, 16#06#),
      2961 => to_slv(opcode_type, 16#B8#),
      2962 => to_slv(opcode_type, 16#0E#),
      2963 => to_slv(opcode_type, 16#06#),
      2964 => to_slv(opcode_type, 16#08#),
      2965 => to_slv(opcode_type, 16#0E#),
      2966 => to_slv(opcode_type, 16#11#),
      2967 => to_slv(opcode_type, 16#05#),
      2968 => to_slv(opcode_type, 16#A5#),
      2969 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#06#),
      2977 => to_slv(opcode_type, 16#06#),
      2978 => to_slv(opcode_type, 16#05#),
      2979 => to_slv(opcode_type, 16#06#),
      2980 => to_slv(opcode_type, 16#0F#),
      2981 => to_slv(opcode_type, 16#0C#),
      2982 => to_slv(opcode_type, 16#06#),
      2983 => to_slv(opcode_type, 16#01#),
      2984 => to_slv(opcode_type, 16#0E#),
      2985 => to_slv(opcode_type, 16#05#),
      2986 => to_slv(opcode_type, 16#0F#),
      2987 => to_slv(opcode_type, 16#07#),
      2988 => to_slv(opcode_type, 16#08#),
      2989 => to_slv(opcode_type, 16#04#),
      2990 => to_slv(opcode_type, 16#0E#),
      2991 => to_slv(opcode_type, 16#08#),
      2992 => to_slv(opcode_type, 16#11#),
      2993 => to_slv(opcode_type, 16#0C#),
      2994 => to_slv(opcode_type, 16#06#),
      2995 => to_slv(opcode_type, 16#07#),
      2996 => to_slv(opcode_type, 16#0B#),
      2997 => to_slv(opcode_type, 16#11#),
      2998 => to_slv(opcode_type, 16#07#),
      2999 => to_slv(opcode_type, 16#0F#),
      3000 => to_slv(opcode_type, 16#0E#),
      3001 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#09#),
      3009 => to_slv(opcode_type, 16#09#),
      3010 => to_slv(opcode_type, 16#06#),
      3011 => to_slv(opcode_type, 16#08#),
      3012 => to_slv(opcode_type, 16#11#),
      3013 => to_slv(opcode_type, 16#0B#),
      3014 => to_slv(opcode_type, 16#06#),
      3015 => to_slv(opcode_type, 16#0E#),
      3016 => to_slv(opcode_type, 16#0E#),
      3017 => to_slv(opcode_type, 16#01#),
      3018 => to_slv(opcode_type, 16#07#),
      3019 => to_slv(opcode_type, 16#0E#),
      3020 => to_slv(opcode_type, 16#0E#),
      3021 => to_slv(opcode_type, 16#09#),
      3022 => to_slv(opcode_type, 16#04#),
      3023 => to_slv(opcode_type, 16#09#),
      3024 => to_slv(opcode_type, 16#E2#),
      3025 => to_slv(opcode_type, 16#B9#),
      3026 => to_slv(opcode_type, 16#07#),
      3027 => to_slv(opcode_type, 16#08#),
      3028 => to_slv(opcode_type, 16#10#),
      3029 => to_slv(opcode_type, 16#0D#),
      3030 => to_slv(opcode_type, 16#08#),
      3031 => to_slv(opcode_type, 16#0F#),
      3032 => to_slv(opcode_type, 16#88#),
      3033 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#09#),
      3041 => to_slv(opcode_type, 16#08#),
      3042 => to_slv(opcode_type, 16#05#),
      3043 => to_slv(opcode_type, 16#03#),
      3044 => to_slv(opcode_type, 16#11#),
      3045 => to_slv(opcode_type, 16#08#),
      3046 => to_slv(opcode_type, 16#03#),
      3047 => to_slv(opcode_type, 16#0B#),
      3048 => to_slv(opcode_type, 16#02#),
      3049 => to_slv(opcode_type, 16#F3#),
      3050 => to_slv(opcode_type, 16#09#),
      3051 => to_slv(opcode_type, 16#09#),
      3052 => to_slv(opcode_type, 16#08#),
      3053 => to_slv(opcode_type, 16#0F#),
      3054 => to_slv(opcode_type, 16#0E#),
      3055 => to_slv(opcode_type, 16#06#),
      3056 => to_slv(opcode_type, 16#0F#),
      3057 => to_slv(opcode_type, 16#0A#),
      3058 => to_slv(opcode_type, 16#07#),
      3059 => to_slv(opcode_type, 16#09#),
      3060 => to_slv(opcode_type, 16#0F#),
      3061 => to_slv(opcode_type, 16#10#),
      3062 => to_slv(opcode_type, 16#09#),
      3063 => to_slv(opcode_type, 16#11#),
      3064 => to_slv(opcode_type, 16#1D#),
      3065 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#08#),
      3073 => to_slv(opcode_type, 16#08#),
      3074 => to_slv(opcode_type, 16#03#),
      3075 => to_slv(opcode_type, 16#04#),
      3076 => to_slv(opcode_type, 16#0C#),
      3077 => to_slv(opcode_type, 16#07#),
      3078 => to_slv(opcode_type, 16#07#),
      3079 => to_slv(opcode_type, 16#10#),
      3080 => to_slv(opcode_type, 16#C0#),
      3081 => to_slv(opcode_type, 16#04#),
      3082 => to_slv(opcode_type, 16#0F#),
      3083 => to_slv(opcode_type, 16#08#),
      3084 => to_slv(opcode_type, 16#08#),
      3085 => to_slv(opcode_type, 16#06#),
      3086 => to_slv(opcode_type, 16#FE#),
      3087 => to_slv(opcode_type, 16#0B#),
      3088 => to_slv(opcode_type, 16#05#),
      3089 => to_slv(opcode_type, 16#0B#),
      3090 => to_slv(opcode_type, 16#08#),
      3091 => to_slv(opcode_type, 16#07#),
      3092 => to_slv(opcode_type, 16#0C#),
      3093 => to_slv(opcode_type, 16#0E#),
      3094 => to_slv(opcode_type, 16#07#),
      3095 => to_slv(opcode_type, 16#0E#),
      3096 => to_slv(opcode_type, 16#61#),
      3097 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#08#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#09#),
      3107 => to_slv(opcode_type, 16#08#),
      3108 => to_slv(opcode_type, 16#63#),
      3109 => to_slv(opcode_type, 16#1C#),
      3110 => to_slv(opcode_type, 16#01#),
      3111 => to_slv(opcode_type, 16#11#),
      3112 => to_slv(opcode_type, 16#09#),
      3113 => to_slv(opcode_type, 16#08#),
      3114 => to_slv(opcode_type, 16#0B#),
      3115 => to_slv(opcode_type, 16#0D#),
      3116 => to_slv(opcode_type, 16#02#),
      3117 => to_slv(opcode_type, 16#10#),
      3118 => to_slv(opcode_type, 16#09#),
      3119 => to_slv(opcode_type, 16#09#),
      3120 => to_slv(opcode_type, 16#03#),
      3121 => to_slv(opcode_type, 16#0D#),
      3122 => to_slv(opcode_type, 16#06#),
      3123 => to_slv(opcode_type, 16#0E#),
      3124 => to_slv(opcode_type, 16#0C#),
      3125 => to_slv(opcode_type, 16#01#),
      3126 => to_slv(opcode_type, 16#07#),
      3127 => to_slv(opcode_type, 16#10#),
      3128 => to_slv(opcode_type, 16#0E#),
      3129 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#08#),
      3137 => to_slv(opcode_type, 16#08#),
      3138 => to_slv(opcode_type, 16#04#),
      3139 => to_slv(opcode_type, 16#09#),
      3140 => to_slv(opcode_type, 16#0C#),
      3141 => to_slv(opcode_type, 16#10#),
      3142 => to_slv(opcode_type, 16#07#),
      3143 => to_slv(opcode_type, 16#07#),
      3144 => to_slv(opcode_type, 16#0E#),
      3145 => to_slv(opcode_type, 16#0E#),
      3146 => to_slv(opcode_type, 16#08#),
      3147 => to_slv(opcode_type, 16#0D#),
      3148 => to_slv(opcode_type, 16#11#),
      3149 => to_slv(opcode_type, 16#06#),
      3150 => to_slv(opcode_type, 16#02#),
      3151 => to_slv(opcode_type, 16#07#),
      3152 => to_slv(opcode_type, 16#0E#),
      3153 => to_slv(opcode_type, 16#11#),
      3154 => to_slv(opcode_type, 16#09#),
      3155 => to_slv(opcode_type, 16#08#),
      3156 => to_slv(opcode_type, 16#11#),
      3157 => to_slv(opcode_type, 16#0E#),
      3158 => to_slv(opcode_type, 16#07#),
      3159 => to_slv(opcode_type, 16#0A#),
      3160 => to_slv(opcode_type, 16#0F#),
      3161 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#09#),
      3169 => to_slv(opcode_type, 16#07#),
      3170 => to_slv(opcode_type, 16#07#),
      3171 => to_slv(opcode_type, 16#06#),
      3172 => to_slv(opcode_type, 16#0F#),
      3173 => to_slv(opcode_type, 16#0D#),
      3174 => to_slv(opcode_type, 16#08#),
      3175 => to_slv(opcode_type, 16#0C#),
      3176 => to_slv(opcode_type, 16#0A#),
      3177 => to_slv(opcode_type, 16#09#),
      3178 => to_slv(opcode_type, 16#07#),
      3179 => to_slv(opcode_type, 16#0F#),
      3180 => to_slv(opcode_type, 16#11#),
      3181 => to_slv(opcode_type, 16#07#),
      3182 => to_slv(opcode_type, 16#0E#),
      3183 => to_slv(opcode_type, 16#32#),
      3184 => to_slv(opcode_type, 16#06#),
      3185 => to_slv(opcode_type, 16#09#),
      3186 => to_slv(opcode_type, 16#04#),
      3187 => to_slv(opcode_type, 16#10#),
      3188 => to_slv(opcode_type, 16#04#),
      3189 => to_slv(opcode_type, 16#11#),
      3190 => to_slv(opcode_type, 16#06#),
      3191 => to_slv(opcode_type, 16#C4#),
      3192 => to_slv(opcode_type, 16#10#),
      3193 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#08#),
      3201 => to_slv(opcode_type, 16#07#),
      3202 => to_slv(opcode_type, 16#03#),
      3203 => to_slv(opcode_type, 16#05#),
      3204 => to_slv(opcode_type, 16#0F#),
      3205 => to_slv(opcode_type, 16#07#),
      3206 => to_slv(opcode_type, 16#08#),
      3207 => to_slv(opcode_type, 16#7A#),
      3208 => to_slv(opcode_type, 16#11#),
      3209 => to_slv(opcode_type, 16#06#),
      3210 => to_slv(opcode_type, 16#0E#),
      3211 => to_slv(opcode_type, 16#11#),
      3212 => to_slv(opcode_type, 16#06#),
      3213 => to_slv(opcode_type, 16#09#),
      3214 => to_slv(opcode_type, 16#07#),
      3215 => to_slv(opcode_type, 16#0C#),
      3216 => to_slv(opcode_type, 16#0B#),
      3217 => to_slv(opcode_type, 16#01#),
      3218 => to_slv(opcode_type, 16#0E#),
      3219 => to_slv(opcode_type, 16#09#),
      3220 => to_slv(opcode_type, 16#05#),
      3221 => to_slv(opcode_type, 16#0A#),
      3222 => to_slv(opcode_type, 16#08#),
      3223 => to_slv(opcode_type, 16#0C#),
      3224 => to_slv(opcode_type, 16#54#),
      3225 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#06#),
      3234 => to_slv(opcode_type, 16#07#),
      3235 => to_slv(opcode_type, 16#02#),
      3236 => to_slv(opcode_type, 16#10#),
      3237 => to_slv(opcode_type, 16#06#),
      3238 => to_slv(opcode_type, 16#0D#),
      3239 => to_slv(opcode_type, 16#11#),
      3240 => to_slv(opcode_type, 16#03#),
      3241 => to_slv(opcode_type, 16#03#),
      3242 => to_slv(opcode_type, 16#0B#),
      3243 => to_slv(opcode_type, 16#09#),
      3244 => to_slv(opcode_type, 16#06#),
      3245 => to_slv(opcode_type, 16#04#),
      3246 => to_slv(opcode_type, 16#0D#),
      3247 => to_slv(opcode_type, 16#07#),
      3248 => to_slv(opcode_type, 16#84#),
      3249 => to_slv(opcode_type, 16#10#),
      3250 => to_slv(opcode_type, 16#06#),
      3251 => to_slv(opcode_type, 16#07#),
      3252 => to_slv(opcode_type, 16#0C#),
      3253 => to_slv(opcode_type, 16#0F#),
      3254 => to_slv(opcode_type, 16#06#),
      3255 => to_slv(opcode_type, 16#0E#),
      3256 => to_slv(opcode_type, 16#0E#),
      3257 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#07#),
      3265 => to_slv(opcode_type, 16#08#),
      3266 => to_slv(opcode_type, 16#01#),
      3267 => to_slv(opcode_type, 16#06#),
      3268 => to_slv(opcode_type, 16#0B#),
      3269 => to_slv(opcode_type, 16#0E#),
      3270 => to_slv(opcode_type, 16#09#),
      3271 => to_slv(opcode_type, 16#03#),
      3272 => to_slv(opcode_type, 16#0F#),
      3273 => to_slv(opcode_type, 16#05#),
      3274 => to_slv(opcode_type, 16#62#),
      3275 => to_slv(opcode_type, 16#08#),
      3276 => to_slv(opcode_type, 16#08#),
      3277 => to_slv(opcode_type, 16#04#),
      3278 => to_slv(opcode_type, 16#0C#),
      3279 => to_slv(opcode_type, 16#09#),
      3280 => to_slv(opcode_type, 16#10#),
      3281 => to_slv(opcode_type, 16#ED#),
      3282 => to_slv(opcode_type, 16#07#),
      3283 => to_slv(opcode_type, 16#08#),
      3284 => to_slv(opcode_type, 16#0C#),
      3285 => to_slv(opcode_type, 16#0F#),
      3286 => to_slv(opcode_type, 16#09#),
      3287 => to_slv(opcode_type, 16#0E#),
      3288 => to_slv(opcode_type, 16#0F#),
      3289 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#06#),
      3297 => to_slv(opcode_type, 16#06#),
      3298 => to_slv(opcode_type, 16#02#),
      3299 => to_slv(opcode_type, 16#03#),
      3300 => to_slv(opcode_type, 16#0B#),
      3301 => to_slv(opcode_type, 16#08#),
      3302 => to_slv(opcode_type, 16#06#),
      3303 => to_slv(opcode_type, 16#11#),
      3304 => to_slv(opcode_type, 16#0B#),
      3305 => to_slv(opcode_type, 16#04#),
      3306 => to_slv(opcode_type, 16#10#),
      3307 => to_slv(opcode_type, 16#09#),
      3308 => to_slv(opcode_type, 16#08#),
      3309 => to_slv(opcode_type, 16#02#),
      3310 => to_slv(opcode_type, 16#74#),
      3311 => to_slv(opcode_type, 16#06#),
      3312 => to_slv(opcode_type, 16#0A#),
      3313 => to_slv(opcode_type, 16#62#),
      3314 => to_slv(opcode_type, 16#08#),
      3315 => to_slv(opcode_type, 16#09#),
      3316 => to_slv(opcode_type, 16#11#),
      3317 => to_slv(opcode_type, 16#11#),
      3318 => to_slv(opcode_type, 16#06#),
      3319 => to_slv(opcode_type, 16#0B#),
      3320 => to_slv(opcode_type, 16#0C#),
      3321 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#07#),
      3329 => to_slv(opcode_type, 16#09#),
      3330 => to_slv(opcode_type, 16#06#),
      3331 => to_slv(opcode_type, 16#04#),
      3332 => to_slv(opcode_type, 16#96#),
      3333 => to_slv(opcode_type, 16#04#),
      3334 => to_slv(opcode_type, 16#0E#),
      3335 => to_slv(opcode_type, 16#09#),
      3336 => to_slv(opcode_type, 16#08#),
      3337 => to_slv(opcode_type, 16#10#),
      3338 => to_slv(opcode_type, 16#0F#),
      3339 => to_slv(opcode_type, 16#06#),
      3340 => to_slv(opcode_type, 16#10#),
      3341 => to_slv(opcode_type, 16#0E#),
      3342 => to_slv(opcode_type, 16#08#),
      3343 => to_slv(opcode_type, 16#06#),
      3344 => to_slv(opcode_type, 16#02#),
      3345 => to_slv(opcode_type, 16#0A#),
      3346 => to_slv(opcode_type, 16#02#),
      3347 => to_slv(opcode_type, 16#10#),
      3348 => to_slv(opcode_type, 16#08#),
      3349 => to_slv(opcode_type, 16#03#),
      3350 => to_slv(opcode_type, 16#0A#),
      3351 => to_slv(opcode_type, 16#02#),
      3352 => to_slv(opcode_type, 16#0C#),
      3353 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#09#),
      3361 => to_slv(opcode_type, 16#06#),
      3362 => to_slv(opcode_type, 16#03#),
      3363 => to_slv(opcode_type, 16#08#),
      3364 => to_slv(opcode_type, 16#0C#),
      3365 => to_slv(opcode_type, 16#10#),
      3366 => to_slv(opcode_type, 16#02#),
      3367 => to_slv(opcode_type, 16#09#),
      3368 => to_slv(opcode_type, 16#0F#),
      3369 => to_slv(opcode_type, 16#0E#),
      3370 => to_slv(opcode_type, 16#06#),
      3371 => to_slv(opcode_type, 16#07#),
      3372 => to_slv(opcode_type, 16#09#),
      3373 => to_slv(opcode_type, 16#0F#),
      3374 => to_slv(opcode_type, 16#0F#),
      3375 => to_slv(opcode_type, 16#09#),
      3376 => to_slv(opcode_type, 16#0F#),
      3377 => to_slv(opcode_type, 16#0C#),
      3378 => to_slv(opcode_type, 16#06#),
      3379 => to_slv(opcode_type, 16#08#),
      3380 => to_slv(opcode_type, 16#11#),
      3381 => to_slv(opcode_type, 16#0B#),
      3382 => to_slv(opcode_type, 16#09#),
      3383 => to_slv(opcode_type, 16#F8#),
      3384 => to_slv(opcode_type, 16#0D#),
      3385 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#09#),
      3393 => to_slv(opcode_type, 16#06#),
      3394 => to_slv(opcode_type, 16#04#),
      3395 => to_slv(opcode_type, 16#01#),
      3396 => to_slv(opcode_type, 16#11#),
      3397 => to_slv(opcode_type, 16#06#),
      3398 => to_slv(opcode_type, 16#06#),
      3399 => to_slv(opcode_type, 16#11#),
      3400 => to_slv(opcode_type, 16#0E#),
      3401 => to_slv(opcode_type, 16#08#),
      3402 => to_slv(opcode_type, 16#10#),
      3403 => to_slv(opcode_type, 16#10#),
      3404 => to_slv(opcode_type, 16#07#),
      3405 => to_slv(opcode_type, 16#07#),
      3406 => to_slv(opcode_type, 16#07#),
      3407 => to_slv(opcode_type, 16#0F#),
      3408 => to_slv(opcode_type, 16#0D#),
      3409 => to_slv(opcode_type, 16#08#),
      3410 => to_slv(opcode_type, 16#0F#),
      3411 => to_slv(opcode_type, 16#0B#),
      3412 => to_slv(opcode_type, 16#06#),
      3413 => to_slv(opcode_type, 16#01#),
      3414 => to_slv(opcode_type, 16#C6#),
      3415 => to_slv(opcode_type, 16#05#),
      3416 => to_slv(opcode_type, 16#0A#),
      3417 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#06#),
      3426 => to_slv(opcode_type, 16#03#),
      3427 => to_slv(opcode_type, 16#09#),
      3428 => to_slv(opcode_type, 16#0B#),
      3429 => to_slv(opcode_type, 16#0C#),
      3430 => to_slv(opcode_type, 16#02#),
      3431 => to_slv(opcode_type, 16#06#),
      3432 => to_slv(opcode_type, 16#0D#),
      3433 => to_slv(opcode_type, 16#0A#),
      3434 => to_slv(opcode_type, 16#09#),
      3435 => to_slv(opcode_type, 16#07#),
      3436 => to_slv(opcode_type, 16#07#),
      3437 => to_slv(opcode_type, 16#0E#),
      3438 => to_slv(opcode_type, 16#0E#),
      3439 => to_slv(opcode_type, 16#06#),
      3440 => to_slv(opcode_type, 16#11#),
      3441 => to_slv(opcode_type, 16#11#),
      3442 => to_slv(opcode_type, 16#09#),
      3443 => to_slv(opcode_type, 16#08#),
      3444 => to_slv(opcode_type, 16#10#),
      3445 => to_slv(opcode_type, 16#11#),
      3446 => to_slv(opcode_type, 16#06#),
      3447 => to_slv(opcode_type, 16#0E#),
      3448 => to_slv(opcode_type, 16#0A#),
      3449 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#06#),
      3457 => to_slv(opcode_type, 16#07#),
      3458 => to_slv(opcode_type, 16#01#),
      3459 => to_slv(opcode_type, 16#01#),
      3460 => to_slv(opcode_type, 16#11#),
      3461 => to_slv(opcode_type, 16#08#),
      3462 => to_slv(opcode_type, 16#05#),
      3463 => to_slv(opcode_type, 16#0B#),
      3464 => to_slv(opcode_type, 16#07#),
      3465 => to_slv(opcode_type, 16#0B#),
      3466 => to_slv(opcode_type, 16#0B#),
      3467 => to_slv(opcode_type, 16#09#),
      3468 => to_slv(opcode_type, 16#08#),
      3469 => to_slv(opcode_type, 16#06#),
      3470 => to_slv(opcode_type, 16#0C#),
      3471 => to_slv(opcode_type, 16#10#),
      3472 => to_slv(opcode_type, 16#07#),
      3473 => to_slv(opcode_type, 16#47#),
      3474 => to_slv(opcode_type, 16#0B#),
      3475 => to_slv(opcode_type, 16#09#),
      3476 => to_slv(opcode_type, 16#06#),
      3477 => to_slv(opcode_type, 16#0C#),
      3478 => to_slv(opcode_type, 16#0A#),
      3479 => to_slv(opcode_type, 16#02#),
      3480 => to_slv(opcode_type, 16#11#),
      3481 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#07#),
      3489 => to_slv(opcode_type, 16#08#),
      3490 => to_slv(opcode_type, 16#06#),
      3491 => to_slv(opcode_type, 16#04#),
      3492 => to_slv(opcode_type, 16#0D#),
      3493 => to_slv(opcode_type, 16#05#),
      3494 => to_slv(opcode_type, 16#0E#),
      3495 => to_slv(opcode_type, 16#06#),
      3496 => to_slv(opcode_type, 16#09#),
      3497 => to_slv(opcode_type, 16#0D#),
      3498 => to_slv(opcode_type, 16#0B#),
      3499 => to_slv(opcode_type, 16#06#),
      3500 => to_slv(opcode_type, 16#0A#),
      3501 => to_slv(opcode_type, 16#0E#),
      3502 => to_slv(opcode_type, 16#06#),
      3503 => to_slv(opcode_type, 16#05#),
      3504 => to_slv(opcode_type, 16#08#),
      3505 => to_slv(opcode_type, 16#10#),
      3506 => to_slv(opcode_type, 16#0D#),
      3507 => to_slv(opcode_type, 16#09#),
      3508 => to_slv(opcode_type, 16#08#),
      3509 => to_slv(opcode_type, 16#11#),
      3510 => to_slv(opcode_type, 16#11#),
      3511 => to_slv(opcode_type, 16#04#),
      3512 => to_slv(opcode_type, 16#0C#),
      3513 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#07#),
      3521 => to_slv(opcode_type, 16#07#),
      3522 => to_slv(opcode_type, 16#06#),
      3523 => to_slv(opcode_type, 16#02#),
      3524 => to_slv(opcode_type, 16#0A#),
      3525 => to_slv(opcode_type, 16#07#),
      3526 => to_slv(opcode_type, 16#10#),
      3527 => to_slv(opcode_type, 16#0D#),
      3528 => to_slv(opcode_type, 16#06#),
      3529 => to_slv(opcode_type, 16#09#),
      3530 => to_slv(opcode_type, 16#11#),
      3531 => to_slv(opcode_type, 16#0A#),
      3532 => to_slv(opcode_type, 16#03#),
      3533 => to_slv(opcode_type, 16#B3#),
      3534 => to_slv(opcode_type, 16#06#),
      3535 => to_slv(opcode_type, 16#09#),
      3536 => to_slv(opcode_type, 16#07#),
      3537 => to_slv(opcode_type, 16#0F#),
      3538 => to_slv(opcode_type, 16#0B#),
      3539 => to_slv(opcode_type, 16#07#),
      3540 => to_slv(opcode_type, 16#0F#),
      3541 => to_slv(opcode_type, 16#0B#),
      3542 => to_slv(opcode_type, 16#04#),
      3543 => to_slv(opcode_type, 16#05#),
      3544 => to_slv(opcode_type, 16#0B#),
      3545 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#09#),
      3553 => to_slv(opcode_type, 16#06#),
      3554 => to_slv(opcode_type, 16#07#),
      3555 => to_slv(opcode_type, 16#08#),
      3556 => to_slv(opcode_type, 16#11#),
      3557 => to_slv(opcode_type, 16#10#),
      3558 => to_slv(opcode_type, 16#06#),
      3559 => to_slv(opcode_type, 16#0A#),
      3560 => to_slv(opcode_type, 16#20#),
      3561 => to_slv(opcode_type, 16#01#),
      3562 => to_slv(opcode_type, 16#03#),
      3563 => to_slv(opcode_type, 16#0A#),
      3564 => to_slv(opcode_type, 16#08#),
      3565 => to_slv(opcode_type, 16#06#),
      3566 => to_slv(opcode_type, 16#02#),
      3567 => to_slv(opcode_type, 16#0D#),
      3568 => to_slv(opcode_type, 16#01#),
      3569 => to_slv(opcode_type, 16#0A#),
      3570 => to_slv(opcode_type, 16#09#),
      3571 => to_slv(opcode_type, 16#06#),
      3572 => to_slv(opcode_type, 16#0E#),
      3573 => to_slv(opcode_type, 16#53#),
      3574 => to_slv(opcode_type, 16#08#),
      3575 => to_slv(opcode_type, 16#0D#),
      3576 => to_slv(opcode_type, 16#10#),
      3577 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#07#),
      3585 => to_slv(opcode_type, 16#06#),
      3586 => to_slv(opcode_type, 16#09#),
      3587 => to_slv(opcode_type, 16#04#),
      3588 => to_slv(opcode_type, 16#11#),
      3589 => to_slv(opcode_type, 16#04#),
      3590 => to_slv(opcode_type, 16#10#),
      3591 => to_slv(opcode_type, 16#01#),
      3592 => to_slv(opcode_type, 16#08#),
      3593 => to_slv(opcode_type, 16#0E#),
      3594 => to_slv(opcode_type, 16#10#),
      3595 => to_slv(opcode_type, 16#06#),
      3596 => to_slv(opcode_type, 16#09#),
      3597 => to_slv(opcode_type, 16#08#),
      3598 => to_slv(opcode_type, 16#0F#),
      3599 => to_slv(opcode_type, 16#0A#),
      3600 => to_slv(opcode_type, 16#03#),
      3601 => to_slv(opcode_type, 16#10#),
      3602 => to_slv(opcode_type, 16#08#),
      3603 => to_slv(opcode_type, 16#06#),
      3604 => to_slv(opcode_type, 16#10#),
      3605 => to_slv(opcode_type, 16#0E#),
      3606 => to_slv(opcode_type, 16#09#),
      3607 => to_slv(opcode_type, 16#10#),
      3608 => to_slv(opcode_type, 16#0D#),
      3609 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#08#),
      3617 => to_slv(opcode_type, 16#06#),
      3618 => to_slv(opcode_type, 16#09#),
      3619 => to_slv(opcode_type, 16#02#),
      3620 => to_slv(opcode_type, 16#0A#),
      3621 => to_slv(opcode_type, 16#05#),
      3622 => to_slv(opcode_type, 16#0D#),
      3623 => to_slv(opcode_type, 16#03#),
      3624 => to_slv(opcode_type, 16#02#),
      3625 => to_slv(opcode_type, 16#10#),
      3626 => to_slv(opcode_type, 16#08#),
      3627 => to_slv(opcode_type, 16#09#),
      3628 => to_slv(opcode_type, 16#08#),
      3629 => to_slv(opcode_type, 16#0A#),
      3630 => to_slv(opcode_type, 16#0B#),
      3631 => to_slv(opcode_type, 16#08#),
      3632 => to_slv(opcode_type, 16#0D#),
      3633 => to_slv(opcode_type, 16#11#),
      3634 => to_slv(opcode_type, 16#06#),
      3635 => to_slv(opcode_type, 16#09#),
      3636 => to_slv(opcode_type, 16#0A#),
      3637 => to_slv(opcode_type, 16#11#),
      3638 => to_slv(opcode_type, 16#09#),
      3639 => to_slv(opcode_type, 16#0B#),
      3640 => to_slv(opcode_type, 16#0D#),
      3641 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#09#),
      3649 => to_slv(opcode_type, 16#06#),
      3650 => to_slv(opcode_type, 16#01#),
      3651 => to_slv(opcode_type, 16#07#),
      3652 => to_slv(opcode_type, 16#0A#),
      3653 => to_slv(opcode_type, 16#BA#),
      3654 => to_slv(opcode_type, 16#06#),
      3655 => to_slv(opcode_type, 16#01#),
      3656 => to_slv(opcode_type, 16#0B#),
      3657 => to_slv(opcode_type, 16#07#),
      3658 => to_slv(opcode_type, 16#0A#),
      3659 => to_slv(opcode_type, 16#11#),
      3660 => to_slv(opcode_type, 16#07#),
      3661 => to_slv(opcode_type, 16#06#),
      3662 => to_slv(opcode_type, 16#09#),
      3663 => to_slv(opcode_type, 16#0B#),
      3664 => to_slv(opcode_type, 16#28#),
      3665 => to_slv(opcode_type, 16#05#),
      3666 => to_slv(opcode_type, 16#0C#),
      3667 => to_slv(opcode_type, 16#07#),
      3668 => to_slv(opcode_type, 16#02#),
      3669 => to_slv(opcode_type, 16#27#),
      3670 => to_slv(opcode_type, 16#09#),
      3671 => to_slv(opcode_type, 16#0B#),
      3672 => to_slv(opcode_type, 16#0A#),
      3673 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#09#),
      3681 => to_slv(opcode_type, 16#08#),
      3682 => to_slv(opcode_type, 16#06#),
      3683 => to_slv(opcode_type, 16#04#),
      3684 => to_slv(opcode_type, 16#0A#),
      3685 => to_slv(opcode_type, 16#02#),
      3686 => to_slv(opcode_type, 16#0B#),
      3687 => to_slv(opcode_type, 16#04#),
      3688 => to_slv(opcode_type, 16#03#),
      3689 => to_slv(opcode_type, 16#0E#),
      3690 => to_slv(opcode_type, 16#07#),
      3691 => to_slv(opcode_type, 16#09#),
      3692 => to_slv(opcode_type, 16#06#),
      3693 => to_slv(opcode_type, 16#0F#),
      3694 => to_slv(opcode_type, 16#0E#),
      3695 => to_slv(opcode_type, 16#07#),
      3696 => to_slv(opcode_type, 16#0C#),
      3697 => to_slv(opcode_type, 16#0C#),
      3698 => to_slv(opcode_type, 16#06#),
      3699 => to_slv(opcode_type, 16#08#),
      3700 => to_slv(opcode_type, 16#0D#),
      3701 => to_slv(opcode_type, 16#0A#),
      3702 => to_slv(opcode_type, 16#06#),
      3703 => to_slv(opcode_type, 16#4E#),
      3704 => to_slv(opcode_type, 16#0A#),
      3705 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#06#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#09#),
      3715 => to_slv(opcode_type, 16#09#),
      3716 => to_slv(opcode_type, 16#0D#),
      3717 => to_slv(opcode_type, 16#21#),
      3718 => to_slv(opcode_type, 16#03#),
      3719 => to_slv(opcode_type, 16#0E#),
      3720 => to_slv(opcode_type, 16#01#),
      3721 => to_slv(opcode_type, 16#04#),
      3722 => to_slv(opcode_type, 16#0C#),
      3723 => to_slv(opcode_type, 16#09#),
      3724 => to_slv(opcode_type, 16#06#),
      3725 => to_slv(opcode_type, 16#05#),
      3726 => to_slv(opcode_type, 16#1A#),
      3727 => to_slv(opcode_type, 16#06#),
      3728 => to_slv(opcode_type, 16#0C#),
      3729 => to_slv(opcode_type, 16#10#),
      3730 => to_slv(opcode_type, 16#08#),
      3731 => to_slv(opcode_type, 16#08#),
      3732 => to_slv(opcode_type, 16#10#),
      3733 => to_slv(opcode_type, 16#E9#),
      3734 => to_slv(opcode_type, 16#06#),
      3735 => to_slv(opcode_type, 16#0D#),
      3736 => to_slv(opcode_type, 16#0C#),
      3737 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#09#),
      3745 => to_slv(opcode_type, 16#09#),
      3746 => to_slv(opcode_type, 16#06#),
      3747 => to_slv(opcode_type, 16#05#),
      3748 => to_slv(opcode_type, 16#0B#),
      3749 => to_slv(opcode_type, 16#04#),
      3750 => to_slv(opcode_type, 16#11#),
      3751 => to_slv(opcode_type, 16#01#),
      3752 => to_slv(opcode_type, 16#07#),
      3753 => to_slv(opcode_type, 16#0D#),
      3754 => to_slv(opcode_type, 16#0E#),
      3755 => to_slv(opcode_type, 16#07#),
      3756 => to_slv(opcode_type, 16#07#),
      3757 => to_slv(opcode_type, 16#01#),
      3758 => to_slv(opcode_type, 16#0A#),
      3759 => to_slv(opcode_type, 16#08#),
      3760 => to_slv(opcode_type, 16#0D#),
      3761 => to_slv(opcode_type, 16#0E#),
      3762 => to_slv(opcode_type, 16#09#),
      3763 => to_slv(opcode_type, 16#09#),
      3764 => to_slv(opcode_type, 16#0F#),
      3765 => to_slv(opcode_type, 16#0D#),
      3766 => to_slv(opcode_type, 16#06#),
      3767 => to_slv(opcode_type, 16#0A#),
      3768 => to_slv(opcode_type, 16#0A#),
      3769 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#09#),
      3777 => to_slv(opcode_type, 16#08#),
      3778 => to_slv(opcode_type, 16#09#),
      3779 => to_slv(opcode_type, 16#02#),
      3780 => to_slv(opcode_type, 16#DF#),
      3781 => to_slv(opcode_type, 16#06#),
      3782 => to_slv(opcode_type, 16#0D#),
      3783 => to_slv(opcode_type, 16#11#),
      3784 => to_slv(opcode_type, 16#03#),
      3785 => to_slv(opcode_type, 16#03#),
      3786 => to_slv(opcode_type, 16#ED#),
      3787 => to_slv(opcode_type, 16#08#),
      3788 => to_slv(opcode_type, 16#09#),
      3789 => to_slv(opcode_type, 16#05#),
      3790 => to_slv(opcode_type, 16#10#),
      3791 => to_slv(opcode_type, 16#09#),
      3792 => to_slv(opcode_type, 16#11#),
      3793 => to_slv(opcode_type, 16#0D#),
      3794 => to_slv(opcode_type, 16#08#),
      3795 => to_slv(opcode_type, 16#06#),
      3796 => to_slv(opcode_type, 16#0D#),
      3797 => to_slv(opcode_type, 16#0E#),
      3798 => to_slv(opcode_type, 16#08#),
      3799 => to_slv(opcode_type, 16#0F#),
      3800 => to_slv(opcode_type, 16#0A#),
      3801 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#09#),
      3809 => to_slv(opcode_type, 16#08#),
      3810 => to_slv(opcode_type, 16#01#),
      3811 => to_slv(opcode_type, 16#07#),
      3812 => to_slv(opcode_type, 16#0B#),
      3813 => to_slv(opcode_type, 16#0F#),
      3814 => to_slv(opcode_type, 16#06#),
      3815 => to_slv(opcode_type, 16#09#),
      3816 => to_slv(opcode_type, 16#0C#),
      3817 => to_slv(opcode_type, 16#0A#),
      3818 => to_slv(opcode_type, 16#05#),
      3819 => to_slv(opcode_type, 16#0B#),
      3820 => to_slv(opcode_type, 16#06#),
      3821 => to_slv(opcode_type, 16#08#),
      3822 => to_slv(opcode_type, 16#02#),
      3823 => to_slv(opcode_type, 16#0E#),
      3824 => to_slv(opcode_type, 16#09#),
      3825 => to_slv(opcode_type, 16#0B#),
      3826 => to_slv(opcode_type, 16#0B#),
      3827 => to_slv(opcode_type, 16#07#),
      3828 => to_slv(opcode_type, 16#06#),
      3829 => to_slv(opcode_type, 16#0D#),
      3830 => to_slv(opcode_type, 16#0D#),
      3831 => to_slv(opcode_type, 16#05#),
      3832 => to_slv(opcode_type, 16#0B#),
      3833 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#08#),
      3841 => to_slv(opcode_type, 16#07#),
      3842 => to_slv(opcode_type, 16#04#),
      3843 => to_slv(opcode_type, 16#02#),
      3844 => to_slv(opcode_type, 16#11#),
      3845 => to_slv(opcode_type, 16#08#),
      3846 => to_slv(opcode_type, 16#06#),
      3847 => to_slv(opcode_type, 16#0F#),
      3848 => to_slv(opcode_type, 16#0B#),
      3849 => to_slv(opcode_type, 16#05#),
      3850 => to_slv(opcode_type, 16#10#),
      3851 => to_slv(opcode_type, 16#06#),
      3852 => to_slv(opcode_type, 16#06#),
      3853 => to_slv(opcode_type, 16#04#),
      3854 => to_slv(opcode_type, 16#0D#),
      3855 => to_slv(opcode_type, 16#08#),
      3856 => to_slv(opcode_type, 16#0A#),
      3857 => to_slv(opcode_type, 16#0C#),
      3858 => to_slv(opcode_type, 16#08#),
      3859 => to_slv(opcode_type, 16#06#),
      3860 => to_slv(opcode_type, 16#11#),
      3861 => to_slv(opcode_type, 16#0C#),
      3862 => to_slv(opcode_type, 16#09#),
      3863 => to_slv(opcode_type, 16#0F#),
      3864 => to_slv(opcode_type, 16#76#),
      3865 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#07#),
      3873 => to_slv(opcode_type, 16#06#),
      3874 => to_slv(opcode_type, 16#02#),
      3875 => to_slv(opcode_type, 16#03#),
      3876 => to_slv(opcode_type, 16#10#),
      3877 => to_slv(opcode_type, 16#07#),
      3878 => to_slv(opcode_type, 16#04#),
      3879 => to_slv(opcode_type, 16#0F#),
      3880 => to_slv(opcode_type, 16#06#),
      3881 => to_slv(opcode_type, 16#0E#),
      3882 => to_slv(opcode_type, 16#10#),
      3883 => to_slv(opcode_type, 16#09#),
      3884 => to_slv(opcode_type, 16#08#),
      3885 => to_slv(opcode_type, 16#02#),
      3886 => to_slv(opcode_type, 16#0A#),
      3887 => to_slv(opcode_type, 16#09#),
      3888 => to_slv(opcode_type, 16#10#),
      3889 => to_slv(opcode_type, 16#0F#),
      3890 => to_slv(opcode_type, 16#08#),
      3891 => to_slv(opcode_type, 16#08#),
      3892 => to_slv(opcode_type, 16#8F#),
      3893 => to_slv(opcode_type, 16#0B#),
      3894 => to_slv(opcode_type, 16#06#),
      3895 => to_slv(opcode_type, 16#92#),
      3896 => to_slv(opcode_type, 16#11#),
      3897 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#08#),
      3905 => to_slv(opcode_type, 16#06#),
      3906 => to_slv(opcode_type, 16#07#),
      3907 => to_slv(opcode_type, 16#09#),
      3908 => to_slv(opcode_type, 16#0E#),
      3909 => to_slv(opcode_type, 16#10#),
      3910 => to_slv(opcode_type, 16#06#),
      3911 => to_slv(opcode_type, 16#0D#),
      3912 => to_slv(opcode_type, 16#11#),
      3913 => to_slv(opcode_type, 16#02#),
      3914 => to_slv(opcode_type, 16#09#),
      3915 => to_slv(opcode_type, 16#68#),
      3916 => to_slv(opcode_type, 16#0D#),
      3917 => to_slv(opcode_type, 16#06#),
      3918 => to_slv(opcode_type, 16#04#),
      3919 => to_slv(opcode_type, 16#09#),
      3920 => to_slv(opcode_type, 16#0A#),
      3921 => to_slv(opcode_type, 16#0A#),
      3922 => to_slv(opcode_type, 16#06#),
      3923 => to_slv(opcode_type, 16#07#),
      3924 => to_slv(opcode_type, 16#0A#),
      3925 => to_slv(opcode_type, 16#0C#),
      3926 => to_slv(opcode_type, 16#06#),
      3927 => to_slv(opcode_type, 16#10#),
      3928 => to_slv(opcode_type, 16#0B#),
      3929 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#08#),
      3937 => to_slv(opcode_type, 16#08#),
      3938 => to_slv(opcode_type, 16#09#),
      3939 => to_slv(opcode_type, 16#06#),
      3940 => to_slv(opcode_type, 16#0C#),
      3941 => to_slv(opcode_type, 16#10#),
      3942 => to_slv(opcode_type, 16#03#),
      3943 => to_slv(opcode_type, 16#0A#),
      3944 => to_slv(opcode_type, 16#08#),
      3945 => to_slv(opcode_type, 16#02#),
      3946 => to_slv(opcode_type, 16#88#),
      3947 => to_slv(opcode_type, 16#08#),
      3948 => to_slv(opcode_type, 16#10#),
      3949 => to_slv(opcode_type, 16#10#),
      3950 => to_slv(opcode_type, 16#07#),
      3951 => to_slv(opcode_type, 16#04#),
      3952 => to_slv(opcode_type, 16#09#),
      3953 => to_slv(opcode_type, 16#CB#),
      3954 => to_slv(opcode_type, 16#10#),
      3955 => to_slv(opcode_type, 16#08#),
      3956 => to_slv(opcode_type, 16#01#),
      3957 => to_slv(opcode_type, 16#0A#),
      3958 => to_slv(opcode_type, 16#09#),
      3959 => to_slv(opcode_type, 16#0B#),
      3960 => to_slv(opcode_type, 16#0F#),
      3961 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#09#),
      3969 => to_slv(opcode_type, 16#06#),
      3970 => to_slv(opcode_type, 16#05#),
      3971 => to_slv(opcode_type, 16#01#),
      3972 => to_slv(opcode_type, 16#26#),
      3973 => to_slv(opcode_type, 16#09#),
      3974 => to_slv(opcode_type, 16#08#),
      3975 => to_slv(opcode_type, 16#0F#),
      3976 => to_slv(opcode_type, 16#0D#),
      3977 => to_slv(opcode_type, 16#06#),
      3978 => to_slv(opcode_type, 16#0D#),
      3979 => to_slv(opcode_type, 16#11#),
      3980 => to_slv(opcode_type, 16#06#),
      3981 => to_slv(opcode_type, 16#07#),
      3982 => to_slv(opcode_type, 16#04#),
      3983 => to_slv(opcode_type, 16#0B#),
      3984 => to_slv(opcode_type, 16#07#),
      3985 => to_slv(opcode_type, 16#0C#),
      3986 => to_slv(opcode_type, 16#0B#),
      3987 => to_slv(opcode_type, 16#07#),
      3988 => to_slv(opcode_type, 16#06#),
      3989 => to_slv(opcode_type, 16#10#),
      3990 => to_slv(opcode_type, 16#0E#),
      3991 => to_slv(opcode_type, 16#02#),
      3992 => to_slv(opcode_type, 16#0C#),
      3993 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#08#),
      4001 => to_slv(opcode_type, 16#06#),
      4002 => to_slv(opcode_type, 16#05#),
      4003 => to_slv(opcode_type, 16#06#),
      4004 => to_slv(opcode_type, 16#0C#),
      4005 => to_slv(opcode_type, 16#0E#),
      4006 => to_slv(opcode_type, 16#02#),
      4007 => to_slv(opcode_type, 16#08#),
      4008 => to_slv(opcode_type, 16#0C#),
      4009 => to_slv(opcode_type, 16#0F#),
      4010 => to_slv(opcode_type, 16#07#),
      4011 => to_slv(opcode_type, 16#09#),
      4012 => to_slv(opcode_type, 16#08#),
      4013 => to_slv(opcode_type, 16#10#),
      4014 => to_slv(opcode_type, 16#0E#),
      4015 => to_slv(opcode_type, 16#07#),
      4016 => to_slv(opcode_type, 16#0D#),
      4017 => to_slv(opcode_type, 16#0B#),
      4018 => to_slv(opcode_type, 16#07#),
      4019 => to_slv(opcode_type, 16#09#),
      4020 => to_slv(opcode_type, 16#33#),
      4021 => to_slv(opcode_type, 16#0C#),
      4022 => to_slv(opcode_type, 16#07#),
      4023 => to_slv(opcode_type, 16#0C#),
      4024 => to_slv(opcode_type, 16#DF#),
      4025 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#07#),
      4033 => to_slv(opcode_type, 16#06#),
      4034 => to_slv(opcode_type, 16#05#),
      4035 => to_slv(opcode_type, 16#06#),
      4036 => to_slv(opcode_type, 16#0C#),
      4037 => to_slv(opcode_type, 16#0A#),
      4038 => to_slv(opcode_type, 16#04#),
      4039 => to_slv(opcode_type, 16#06#),
      4040 => to_slv(opcode_type, 16#B0#),
      4041 => to_slv(opcode_type, 16#7C#),
      4042 => to_slv(opcode_type, 16#07#),
      4043 => to_slv(opcode_type, 16#07#),
      4044 => to_slv(opcode_type, 16#06#),
      4045 => to_slv(opcode_type, 16#5D#),
      4046 => to_slv(opcode_type, 16#0F#),
      4047 => to_slv(opcode_type, 16#07#),
      4048 => to_slv(opcode_type, 16#0A#),
      4049 => to_slv(opcode_type, 16#0F#),
      4050 => to_slv(opcode_type, 16#07#),
      4051 => to_slv(opcode_type, 16#06#),
      4052 => to_slv(opcode_type, 16#0E#),
      4053 => to_slv(opcode_type, 16#0A#),
      4054 => to_slv(opcode_type, 16#07#),
      4055 => to_slv(opcode_type, 16#20#),
      4056 => to_slv(opcode_type, 16#11#),
      4057 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#08#),
      4066 => to_slv(opcode_type, 16#01#),
      4067 => to_slv(opcode_type, 16#04#),
      4068 => to_slv(opcode_type, 16#10#),
      4069 => to_slv(opcode_type, 16#08#),
      4070 => to_slv(opcode_type, 16#09#),
      4071 => to_slv(opcode_type, 16#17#),
      4072 => to_slv(opcode_type, 16#0D#),
      4073 => to_slv(opcode_type, 16#08#),
      4074 => to_slv(opcode_type, 16#0D#),
      4075 => to_slv(opcode_type, 16#11#),
      4076 => to_slv(opcode_type, 16#06#),
      4077 => to_slv(opcode_type, 16#08#),
      4078 => to_slv(opcode_type, 16#06#),
      4079 => to_slv(opcode_type, 16#10#),
      4080 => to_slv(opcode_type, 16#0A#),
      4081 => to_slv(opcode_type, 16#02#),
      4082 => to_slv(opcode_type, 16#0D#),
      4083 => to_slv(opcode_type, 16#07#),
      4084 => to_slv(opcode_type, 16#09#),
      4085 => to_slv(opcode_type, 16#11#),
      4086 => to_slv(opcode_type, 16#0D#),
      4087 => to_slv(opcode_type, 16#05#),
      4088 => to_slv(opcode_type, 16#0E#),
      4089 to 4095 => (others => '0')
  ),

    -- Bin `26`...
    25 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#08#),
      1 => to_slv(opcode_type, 16#09#),
      2 => to_slv(opcode_type, 16#02#),
      3 => to_slv(opcode_type, 16#04#),
      4 => to_slv(opcode_type, 16#0B#),
      5 => to_slv(opcode_type, 16#09#),
      6 => to_slv(opcode_type, 16#01#),
      7 => to_slv(opcode_type, 16#0E#),
      8 => to_slv(opcode_type, 16#07#),
      9 => to_slv(opcode_type, 16#0D#),
      10 => to_slv(opcode_type, 16#0B#),
      11 => to_slv(opcode_type, 16#07#),
      12 => to_slv(opcode_type, 16#08#),
      13 => to_slv(opcode_type, 16#08#),
      14 => to_slv(opcode_type, 16#64#),
      15 => to_slv(opcode_type, 16#10#),
      16 => to_slv(opcode_type, 16#07#),
      17 => to_slv(opcode_type, 16#0B#),
      18 => to_slv(opcode_type, 16#10#),
      19 => to_slv(opcode_type, 16#09#),
      20 => to_slv(opcode_type, 16#06#),
      21 => to_slv(opcode_type, 16#0C#),
      22 => to_slv(opcode_type, 16#0F#),
      23 => to_slv(opcode_type, 16#06#),
      24 => to_slv(opcode_type, 16#10#),
      25 => to_slv(opcode_type, 16#0B#),
      26 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#09#),
      33 => to_slv(opcode_type, 16#07#),
      34 => to_slv(opcode_type, 16#08#),
      35 => to_slv(opcode_type, 16#04#),
      36 => to_slv(opcode_type, 16#0B#),
      37 => to_slv(opcode_type, 16#04#),
      38 => to_slv(opcode_type, 16#0C#),
      39 => to_slv(opcode_type, 16#08#),
      40 => to_slv(opcode_type, 16#03#),
      41 => to_slv(opcode_type, 16#0D#),
      42 => to_slv(opcode_type, 16#02#),
      43 => to_slv(opcode_type, 16#0D#),
      44 => to_slv(opcode_type, 16#07#),
      45 => to_slv(opcode_type, 16#07#),
      46 => to_slv(opcode_type, 16#07#),
      47 => to_slv(opcode_type, 16#0C#),
      48 => to_slv(opcode_type, 16#0F#),
      49 => to_slv(opcode_type, 16#03#),
      50 => to_slv(opcode_type, 16#0C#),
      51 => to_slv(opcode_type, 16#09#),
      52 => to_slv(opcode_type, 16#07#),
      53 => to_slv(opcode_type, 16#0B#),
      54 => to_slv(opcode_type, 16#0E#),
      55 => to_slv(opcode_type, 16#07#),
      56 => to_slv(opcode_type, 16#0F#),
      57 => to_slv(opcode_type, 16#0F#),
      58 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#09#),
      65 => to_slv(opcode_type, 16#09#),
      66 => to_slv(opcode_type, 16#02#),
      67 => to_slv(opcode_type, 16#08#),
      68 => to_slv(opcode_type, 16#10#),
      69 => to_slv(opcode_type, 16#0F#),
      70 => to_slv(opcode_type, 16#09#),
      71 => to_slv(opcode_type, 16#08#),
      72 => to_slv(opcode_type, 16#11#),
      73 => to_slv(opcode_type, 16#0D#),
      74 => to_slv(opcode_type, 16#03#),
      75 => to_slv(opcode_type, 16#0A#),
      76 => to_slv(opcode_type, 16#09#),
      77 => to_slv(opcode_type, 16#09#),
      78 => to_slv(opcode_type, 16#07#),
      79 => to_slv(opcode_type, 16#0D#),
      80 => to_slv(opcode_type, 16#0B#),
      81 => to_slv(opcode_type, 16#07#),
      82 => to_slv(opcode_type, 16#0F#),
      83 => to_slv(opcode_type, 16#0E#),
      84 => to_slv(opcode_type, 16#07#),
      85 => to_slv(opcode_type, 16#01#),
      86 => to_slv(opcode_type, 16#11#),
      87 => to_slv(opcode_type, 16#06#),
      88 => to_slv(opcode_type, 16#0A#),
      89 => to_slv(opcode_type, 16#0C#),
      90 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#07#),
      97 => to_slv(opcode_type, 16#06#),
      98 => to_slv(opcode_type, 16#09#),
      99 => to_slv(opcode_type, 16#06#),
      100 => to_slv(opcode_type, 16#0F#),
      101 => to_slv(opcode_type, 16#9E#),
      102 => to_slv(opcode_type, 16#04#),
      103 => to_slv(opcode_type, 16#10#),
      104 => to_slv(opcode_type, 16#06#),
      105 => to_slv(opcode_type, 16#02#),
      106 => to_slv(opcode_type, 16#0D#),
      107 => to_slv(opcode_type, 16#03#),
      108 => to_slv(opcode_type, 16#0F#),
      109 => to_slv(opcode_type, 16#08#),
      110 => to_slv(opcode_type, 16#09#),
      111 => to_slv(opcode_type, 16#04#),
      112 => to_slv(opcode_type, 16#0D#),
      113 => to_slv(opcode_type, 16#05#),
      114 => to_slv(opcode_type, 16#0F#),
      115 => to_slv(opcode_type, 16#06#),
      116 => to_slv(opcode_type, 16#08#),
      117 => to_slv(opcode_type, 16#0F#),
      118 => to_slv(opcode_type, 16#10#),
      119 => to_slv(opcode_type, 16#08#),
      120 => to_slv(opcode_type, 16#0A#),
      121 => to_slv(opcode_type, 16#0F#),
      122 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#08#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#03#),
      131 => to_slv(opcode_type, 16#09#),
      132 => to_slv(opcode_type, 16#0D#),
      133 => to_slv(opcode_type, 16#E1#),
      134 => to_slv(opcode_type, 16#08#),
      135 => to_slv(opcode_type, 16#01#),
      136 => to_slv(opcode_type, 16#0A#),
      137 => to_slv(opcode_type, 16#08#),
      138 => to_slv(opcode_type, 16#65#),
      139 => to_slv(opcode_type, 16#10#),
      140 => to_slv(opcode_type, 16#09#),
      141 => to_slv(opcode_type, 16#08#),
      142 => to_slv(opcode_type, 16#02#),
      143 => to_slv(opcode_type, 16#0A#),
      144 => to_slv(opcode_type, 16#07#),
      145 => to_slv(opcode_type, 16#0F#),
      146 => to_slv(opcode_type, 16#2B#),
      147 => to_slv(opcode_type, 16#09#),
      148 => to_slv(opcode_type, 16#09#),
      149 => to_slv(opcode_type, 16#0C#),
      150 => to_slv(opcode_type, 16#B7#),
      151 => to_slv(opcode_type, 16#07#),
      152 => to_slv(opcode_type, 16#0A#),
      153 => to_slv(opcode_type, 16#11#),
      154 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#09#),
      161 => to_slv(opcode_type, 16#06#),
      162 => to_slv(opcode_type, 16#08#),
      163 => to_slv(opcode_type, 16#03#),
      164 => to_slv(opcode_type, 16#0C#),
      165 => to_slv(opcode_type, 16#06#),
      166 => to_slv(opcode_type, 16#10#),
      167 => to_slv(opcode_type, 16#0E#),
      168 => to_slv(opcode_type, 16#03#),
      169 => to_slv(opcode_type, 16#09#),
      170 => to_slv(opcode_type, 16#0D#),
      171 => to_slv(opcode_type, 16#0E#),
      172 => to_slv(opcode_type, 16#07#),
      173 => to_slv(opcode_type, 16#08#),
      174 => to_slv(opcode_type, 16#07#),
      175 => to_slv(opcode_type, 16#0C#),
      176 => to_slv(opcode_type, 16#0A#),
      177 => to_slv(opcode_type, 16#01#),
      178 => to_slv(opcode_type, 16#0A#),
      179 => to_slv(opcode_type, 16#07#),
      180 => to_slv(opcode_type, 16#07#),
      181 => to_slv(opcode_type, 16#0B#),
      182 => to_slv(opcode_type, 16#0F#),
      183 => to_slv(opcode_type, 16#08#),
      184 => to_slv(opcode_type, 16#D6#),
      185 => to_slv(opcode_type, 16#0A#),
      186 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#06#),
      193 => to_slv(opcode_type, 16#09#),
      194 => to_slv(opcode_type, 16#04#),
      195 => to_slv(opcode_type, 16#08#),
      196 => to_slv(opcode_type, 16#0D#),
      197 => to_slv(opcode_type, 16#A6#),
      198 => to_slv(opcode_type, 16#06#),
      199 => to_slv(opcode_type, 16#07#),
      200 => to_slv(opcode_type, 16#0F#),
      201 => to_slv(opcode_type, 16#0C#),
      202 => to_slv(opcode_type, 16#04#),
      203 => to_slv(opcode_type, 16#10#),
      204 => to_slv(opcode_type, 16#09#),
      205 => to_slv(opcode_type, 16#06#),
      206 => to_slv(opcode_type, 16#04#),
      207 => to_slv(opcode_type, 16#0C#),
      208 => to_slv(opcode_type, 16#08#),
      209 => to_slv(opcode_type, 16#0E#),
      210 => to_slv(opcode_type, 16#0B#),
      211 => to_slv(opcode_type, 16#06#),
      212 => to_slv(opcode_type, 16#06#),
      213 => to_slv(opcode_type, 16#0E#),
      214 => to_slv(opcode_type, 16#0D#),
      215 => to_slv(opcode_type, 16#09#),
      216 => to_slv(opcode_type, 16#11#),
      217 => to_slv(opcode_type, 16#0D#),
      218 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#09#),
      225 => to_slv(opcode_type, 16#06#),
      226 => to_slv(opcode_type, 16#01#),
      227 => to_slv(opcode_type, 16#02#),
      228 => to_slv(opcode_type, 16#11#),
      229 => to_slv(opcode_type, 16#06#),
      230 => to_slv(opcode_type, 16#03#),
      231 => to_slv(opcode_type, 16#0C#),
      232 => to_slv(opcode_type, 16#07#),
      233 => to_slv(opcode_type, 16#10#),
      234 => to_slv(opcode_type, 16#10#),
      235 => to_slv(opcode_type, 16#07#),
      236 => to_slv(opcode_type, 16#06#),
      237 => to_slv(opcode_type, 16#09#),
      238 => to_slv(opcode_type, 16#0E#),
      239 => to_slv(opcode_type, 16#0F#),
      240 => to_slv(opcode_type, 16#08#),
      241 => to_slv(opcode_type, 16#0A#),
      242 => to_slv(opcode_type, 16#11#),
      243 => to_slv(opcode_type, 16#09#),
      244 => to_slv(opcode_type, 16#08#),
      245 => to_slv(opcode_type, 16#FE#),
      246 => to_slv(opcode_type, 16#11#),
      247 => to_slv(opcode_type, 16#07#),
      248 => to_slv(opcode_type, 16#10#),
      249 => to_slv(opcode_type, 16#10#),
      250 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#08#),
      257 => to_slv(opcode_type, 16#08#),
      258 => to_slv(opcode_type, 16#01#),
      259 => to_slv(opcode_type, 16#01#),
      260 => to_slv(opcode_type, 16#0F#),
      261 => to_slv(opcode_type, 16#08#),
      262 => to_slv(opcode_type, 16#01#),
      263 => to_slv(opcode_type, 16#0B#),
      264 => to_slv(opcode_type, 16#07#),
      265 => to_slv(opcode_type, 16#0F#),
      266 => to_slv(opcode_type, 16#0C#),
      267 => to_slv(opcode_type, 16#07#),
      268 => to_slv(opcode_type, 16#06#),
      269 => to_slv(opcode_type, 16#07#),
      270 => to_slv(opcode_type, 16#0E#),
      271 => to_slv(opcode_type, 16#0F#),
      272 => to_slv(opcode_type, 16#09#),
      273 => to_slv(opcode_type, 16#11#),
      274 => to_slv(opcode_type, 16#E9#),
      275 => to_slv(opcode_type, 16#09#),
      276 => to_slv(opcode_type, 16#09#),
      277 => to_slv(opcode_type, 16#10#),
      278 => to_slv(opcode_type, 16#0F#),
      279 => to_slv(opcode_type, 16#07#),
      280 => to_slv(opcode_type, 16#0E#),
      281 => to_slv(opcode_type, 16#2A#),
      282 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#06#),
      289 => to_slv(opcode_type, 16#07#),
      290 => to_slv(opcode_type, 16#04#),
      291 => to_slv(opcode_type, 16#03#),
      292 => to_slv(opcode_type, 16#0D#),
      293 => to_slv(opcode_type, 16#08#),
      294 => to_slv(opcode_type, 16#01#),
      295 => to_slv(opcode_type, 16#0F#),
      296 => to_slv(opcode_type, 16#09#),
      297 => to_slv(opcode_type, 16#0F#),
      298 => to_slv(opcode_type, 16#10#),
      299 => to_slv(opcode_type, 16#09#),
      300 => to_slv(opcode_type, 16#06#),
      301 => to_slv(opcode_type, 16#07#),
      302 => to_slv(opcode_type, 16#0B#),
      303 => to_slv(opcode_type, 16#0E#),
      304 => to_slv(opcode_type, 16#07#),
      305 => to_slv(opcode_type, 16#C3#),
      306 => to_slv(opcode_type, 16#0B#),
      307 => to_slv(opcode_type, 16#08#),
      308 => to_slv(opcode_type, 16#09#),
      309 => to_slv(opcode_type, 16#21#),
      310 => to_slv(opcode_type, 16#0B#),
      311 => to_slv(opcode_type, 16#06#),
      312 => to_slv(opcode_type, 16#0D#),
      313 => to_slv(opcode_type, 16#11#),
      314 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#09#),
      321 => to_slv(opcode_type, 16#08#),
      322 => to_slv(opcode_type, 16#09#),
      323 => to_slv(opcode_type, 16#07#),
      324 => to_slv(opcode_type, 16#0B#),
      325 => to_slv(opcode_type, 16#0E#),
      326 => to_slv(opcode_type, 16#08#),
      327 => to_slv(opcode_type, 16#0C#),
      328 => to_slv(opcode_type, 16#0E#),
      329 => to_slv(opcode_type, 16#04#),
      330 => to_slv(opcode_type, 16#06#),
      331 => to_slv(opcode_type, 16#0D#),
      332 => to_slv(opcode_type, 16#0F#),
      333 => to_slv(opcode_type, 16#07#),
      334 => to_slv(opcode_type, 16#08#),
      335 => to_slv(opcode_type, 16#02#),
      336 => to_slv(opcode_type, 16#0F#),
      337 => to_slv(opcode_type, 16#09#),
      338 => to_slv(opcode_type, 16#0F#),
      339 => to_slv(opcode_type, 16#0F#),
      340 => to_slv(opcode_type, 16#09#),
      341 => to_slv(opcode_type, 16#04#),
      342 => to_slv(opcode_type, 16#0E#),
      343 => to_slv(opcode_type, 16#07#),
      344 => to_slv(opcode_type, 16#0B#),
      345 => to_slv(opcode_type, 16#0A#),
      346 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#08#),
      353 => to_slv(opcode_type, 16#07#),
      354 => to_slv(opcode_type, 16#07#),
      355 => to_slv(opcode_type, 16#04#),
      356 => to_slv(opcode_type, 16#0B#),
      357 => to_slv(opcode_type, 16#04#),
      358 => to_slv(opcode_type, 16#0B#),
      359 => to_slv(opcode_type, 16#04#),
      360 => to_slv(opcode_type, 16#08#),
      361 => to_slv(opcode_type, 16#0C#),
      362 => to_slv(opcode_type, 16#10#),
      363 => to_slv(opcode_type, 16#06#),
      364 => to_slv(opcode_type, 16#07#),
      365 => to_slv(opcode_type, 16#07#),
      366 => to_slv(opcode_type, 16#DB#),
      367 => to_slv(opcode_type, 16#D0#),
      368 => to_slv(opcode_type, 16#08#),
      369 => to_slv(opcode_type, 16#11#),
      370 => to_slv(opcode_type, 16#98#),
      371 => to_slv(opcode_type, 16#06#),
      372 => to_slv(opcode_type, 16#07#),
      373 => to_slv(opcode_type, 16#0B#),
      374 => to_slv(opcode_type, 16#0C#),
      375 => to_slv(opcode_type, 16#06#),
      376 => to_slv(opcode_type, 16#0E#),
      377 => to_slv(opcode_type, 16#0E#),
      378 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#07#),
      385 => to_slv(opcode_type, 16#07#),
      386 => to_slv(opcode_type, 16#01#),
      387 => to_slv(opcode_type, 16#07#),
      388 => to_slv(opcode_type, 16#11#),
      389 => to_slv(opcode_type, 16#0A#),
      390 => to_slv(opcode_type, 16#08#),
      391 => to_slv(opcode_type, 16#05#),
      392 => to_slv(opcode_type, 16#0B#),
      393 => to_slv(opcode_type, 16#07#),
      394 => to_slv(opcode_type, 16#0A#),
      395 => to_slv(opcode_type, 16#0C#),
      396 => to_slv(opcode_type, 16#08#),
      397 => to_slv(opcode_type, 16#09#),
      398 => to_slv(opcode_type, 16#06#),
      399 => to_slv(opcode_type, 16#0A#),
      400 => to_slv(opcode_type, 16#0D#),
      401 => to_slv(opcode_type, 16#04#),
      402 => to_slv(opcode_type, 16#EA#),
      403 => to_slv(opcode_type, 16#07#),
      404 => to_slv(opcode_type, 16#08#),
      405 => to_slv(opcode_type, 16#0E#),
      406 => to_slv(opcode_type, 16#10#),
      407 => to_slv(opcode_type, 16#09#),
      408 => to_slv(opcode_type, 16#0D#),
      409 => to_slv(opcode_type, 16#0A#),
      410 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#07#),
      417 => to_slv(opcode_type, 16#06#),
      418 => to_slv(opcode_type, 16#07#),
      419 => to_slv(opcode_type, 16#07#),
      420 => to_slv(opcode_type, 16#0B#),
      421 => to_slv(opcode_type, 16#0F#),
      422 => to_slv(opcode_type, 16#07#),
      423 => to_slv(opcode_type, 16#0E#),
      424 => to_slv(opcode_type, 16#0D#),
      425 => to_slv(opcode_type, 16#07#),
      426 => to_slv(opcode_type, 16#09#),
      427 => to_slv(opcode_type, 16#0C#),
      428 => to_slv(opcode_type, 16#0E#),
      429 => to_slv(opcode_type, 16#07#),
      430 => to_slv(opcode_type, 16#0F#),
      431 => to_slv(opcode_type, 16#0D#),
      432 => to_slv(opcode_type, 16#06#),
      433 => to_slv(opcode_type, 16#01#),
      434 => to_slv(opcode_type, 16#01#),
      435 => to_slv(opcode_type, 16#0A#),
      436 => to_slv(opcode_type, 16#08#),
      437 => to_slv(opcode_type, 16#08#),
      438 => to_slv(opcode_type, 16#0F#),
      439 => to_slv(opcode_type, 16#0B#),
      440 => to_slv(opcode_type, 16#04#),
      441 => to_slv(opcode_type, 16#EB#),
      442 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#06#),
      449 => to_slv(opcode_type, 16#07#),
      450 => to_slv(opcode_type, 16#07#),
      451 => to_slv(opcode_type, 16#07#),
      452 => to_slv(opcode_type, 16#0F#),
      453 => to_slv(opcode_type, 16#0C#),
      454 => to_slv(opcode_type, 16#01#),
      455 => to_slv(opcode_type, 16#10#),
      456 => to_slv(opcode_type, 16#05#),
      457 => to_slv(opcode_type, 16#05#),
      458 => to_slv(opcode_type, 16#0F#),
      459 => to_slv(opcode_type, 16#07#),
      460 => to_slv(opcode_type, 16#06#),
      461 => to_slv(opcode_type, 16#07#),
      462 => to_slv(opcode_type, 16#0D#),
      463 => to_slv(opcode_type, 16#10#),
      464 => to_slv(opcode_type, 16#08#),
      465 => to_slv(opcode_type, 16#0F#),
      466 => to_slv(opcode_type, 16#11#),
      467 => to_slv(opcode_type, 16#08#),
      468 => to_slv(opcode_type, 16#06#),
      469 => to_slv(opcode_type, 16#0C#),
      470 => to_slv(opcode_type, 16#1F#),
      471 => to_slv(opcode_type, 16#09#),
      472 => to_slv(opcode_type, 16#0E#),
      473 => to_slv(opcode_type, 16#0D#),
      474 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#07#),
      481 => to_slv(opcode_type, 16#09#),
      482 => to_slv(opcode_type, 16#09#),
      483 => to_slv(opcode_type, 16#06#),
      484 => to_slv(opcode_type, 16#0D#),
      485 => to_slv(opcode_type, 16#0D#),
      486 => to_slv(opcode_type, 16#01#),
      487 => to_slv(opcode_type, 16#0E#),
      488 => to_slv(opcode_type, 16#01#),
      489 => to_slv(opcode_type, 16#09#),
      490 => to_slv(opcode_type, 16#0E#),
      491 => to_slv(opcode_type, 16#0B#),
      492 => to_slv(opcode_type, 16#09#),
      493 => to_slv(opcode_type, 16#06#),
      494 => to_slv(opcode_type, 16#04#),
      495 => to_slv(opcode_type, 16#4E#),
      496 => to_slv(opcode_type, 16#06#),
      497 => to_slv(opcode_type, 16#10#),
      498 => to_slv(opcode_type, 16#0B#),
      499 => to_slv(opcode_type, 16#06#),
      500 => to_slv(opcode_type, 16#07#),
      501 => to_slv(opcode_type, 16#11#),
      502 => to_slv(opcode_type, 16#ED#),
      503 => to_slv(opcode_type, 16#09#),
      504 => to_slv(opcode_type, 16#BB#),
      505 => to_slv(opcode_type, 16#0C#),
      506 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#07#),
      513 => to_slv(opcode_type, 16#07#),
      514 => to_slv(opcode_type, 16#04#),
      515 => to_slv(opcode_type, 16#01#),
      516 => to_slv(opcode_type, 16#0D#),
      517 => to_slv(opcode_type, 16#09#),
      518 => to_slv(opcode_type, 16#09#),
      519 => to_slv(opcode_type, 16#0F#),
      520 => to_slv(opcode_type, 16#0D#),
      521 => to_slv(opcode_type, 16#03#),
      522 => to_slv(opcode_type, 16#0A#),
      523 => to_slv(opcode_type, 16#09#),
      524 => to_slv(opcode_type, 16#07#),
      525 => to_slv(opcode_type, 16#09#),
      526 => to_slv(opcode_type, 16#10#),
      527 => to_slv(opcode_type, 16#10#),
      528 => to_slv(opcode_type, 16#06#),
      529 => to_slv(opcode_type, 16#0E#),
      530 => to_slv(opcode_type, 16#0C#),
      531 => to_slv(opcode_type, 16#07#),
      532 => to_slv(opcode_type, 16#08#),
      533 => to_slv(opcode_type, 16#ED#),
      534 => to_slv(opcode_type, 16#11#),
      535 => to_slv(opcode_type, 16#06#),
      536 => to_slv(opcode_type, 16#11#),
      537 => to_slv(opcode_type, 16#11#),
      538 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#06#),
      545 => to_slv(opcode_type, 16#06#),
      546 => to_slv(opcode_type, 16#07#),
      547 => to_slv(opcode_type, 16#04#),
      548 => to_slv(opcode_type, 16#9D#),
      549 => to_slv(opcode_type, 16#07#),
      550 => to_slv(opcode_type, 16#0E#),
      551 => to_slv(opcode_type, 16#0D#),
      552 => to_slv(opcode_type, 16#05#),
      553 => to_slv(opcode_type, 16#01#),
      554 => to_slv(opcode_type, 16#0F#),
      555 => to_slv(opcode_type, 16#06#),
      556 => to_slv(opcode_type, 16#09#),
      557 => to_slv(opcode_type, 16#07#),
      558 => to_slv(opcode_type, 16#0D#),
      559 => to_slv(opcode_type, 16#10#),
      560 => to_slv(opcode_type, 16#09#),
      561 => to_slv(opcode_type, 16#0A#),
      562 => to_slv(opcode_type, 16#11#),
      563 => to_slv(opcode_type, 16#06#),
      564 => to_slv(opcode_type, 16#07#),
      565 => to_slv(opcode_type, 16#0C#),
      566 => to_slv(opcode_type, 16#0D#),
      567 => to_slv(opcode_type, 16#09#),
      568 => to_slv(opcode_type, 16#10#),
      569 => to_slv(opcode_type, 16#0C#),
      570 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#06#),
      577 => to_slv(opcode_type, 16#09#),
      578 => to_slv(opcode_type, 16#03#),
      579 => to_slv(opcode_type, 16#09#),
      580 => to_slv(opcode_type, 16#0A#),
      581 => to_slv(opcode_type, 16#0F#),
      582 => to_slv(opcode_type, 16#06#),
      583 => to_slv(opcode_type, 16#09#),
      584 => to_slv(opcode_type, 16#95#),
      585 => to_slv(opcode_type, 16#10#),
      586 => to_slv(opcode_type, 16#06#),
      587 => to_slv(opcode_type, 16#10#),
      588 => to_slv(opcode_type, 16#0E#),
      589 => to_slv(opcode_type, 16#09#),
      590 => to_slv(opcode_type, 16#06#),
      591 => to_slv(opcode_type, 16#07#),
      592 => to_slv(opcode_type, 16#65#),
      593 => to_slv(opcode_type, 16#10#),
      594 => to_slv(opcode_type, 16#09#),
      595 => to_slv(opcode_type, 16#0D#),
      596 => to_slv(opcode_type, 16#0D#),
      597 => to_slv(opcode_type, 16#07#),
      598 => to_slv(opcode_type, 16#07#),
      599 => to_slv(opcode_type, 16#0E#),
      600 => to_slv(opcode_type, 16#0A#),
      601 => to_slv(opcode_type, 16#0E#),
      602 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#09#),
      609 => to_slv(opcode_type, 16#08#),
      610 => to_slv(opcode_type, 16#02#),
      611 => to_slv(opcode_type, 16#08#),
      612 => to_slv(opcode_type, 16#F6#),
      613 => to_slv(opcode_type, 16#0F#),
      614 => to_slv(opcode_type, 16#07#),
      615 => to_slv(opcode_type, 16#01#),
      616 => to_slv(opcode_type, 16#0E#),
      617 => to_slv(opcode_type, 16#05#),
      618 => to_slv(opcode_type, 16#0B#),
      619 => to_slv(opcode_type, 16#09#),
      620 => to_slv(opcode_type, 16#09#),
      621 => to_slv(opcode_type, 16#09#),
      622 => to_slv(opcode_type, 16#0C#),
      623 => to_slv(opcode_type, 16#BB#),
      624 => to_slv(opcode_type, 16#07#),
      625 => to_slv(opcode_type, 16#E1#),
      626 => to_slv(opcode_type, 16#0A#),
      627 => to_slv(opcode_type, 16#08#),
      628 => to_slv(opcode_type, 16#09#),
      629 => to_slv(opcode_type, 16#0E#),
      630 => to_slv(opcode_type, 16#0C#),
      631 => to_slv(opcode_type, 16#07#),
      632 => to_slv(opcode_type, 16#10#),
      633 => to_slv(opcode_type, 16#10#),
      634 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#09#),
      641 => to_slv(opcode_type, 16#08#),
      642 => to_slv(opcode_type, 16#01#),
      643 => to_slv(opcode_type, 16#03#),
      644 => to_slv(opcode_type, 16#0C#),
      645 => to_slv(opcode_type, 16#07#),
      646 => to_slv(opcode_type, 16#06#),
      647 => to_slv(opcode_type, 16#0E#),
      648 => to_slv(opcode_type, 16#0C#),
      649 => to_slv(opcode_type, 16#07#),
      650 => to_slv(opcode_type, 16#0C#),
      651 => to_slv(opcode_type, 16#0F#),
      652 => to_slv(opcode_type, 16#07#),
      653 => to_slv(opcode_type, 16#07#),
      654 => to_slv(opcode_type, 16#02#),
      655 => to_slv(opcode_type, 16#0B#),
      656 => to_slv(opcode_type, 16#06#),
      657 => to_slv(opcode_type, 16#0F#),
      658 => to_slv(opcode_type, 16#0A#),
      659 => to_slv(opcode_type, 16#08#),
      660 => to_slv(opcode_type, 16#06#),
      661 => to_slv(opcode_type, 16#10#),
      662 => to_slv(opcode_type, 16#0B#),
      663 => to_slv(opcode_type, 16#08#),
      664 => to_slv(opcode_type, 16#11#),
      665 => to_slv(opcode_type, 16#0E#),
      666 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#06#),
      673 => to_slv(opcode_type, 16#07#),
      674 => to_slv(opcode_type, 16#04#),
      675 => to_slv(opcode_type, 16#03#),
      676 => to_slv(opcode_type, 16#11#),
      677 => to_slv(opcode_type, 16#08#),
      678 => to_slv(opcode_type, 16#08#),
      679 => to_slv(opcode_type, 16#23#),
      680 => to_slv(opcode_type, 16#0F#),
      681 => to_slv(opcode_type, 16#02#),
      682 => to_slv(opcode_type, 16#11#),
      683 => to_slv(opcode_type, 16#07#),
      684 => to_slv(opcode_type, 16#09#),
      685 => to_slv(opcode_type, 16#09#),
      686 => to_slv(opcode_type, 16#0D#),
      687 => to_slv(opcode_type, 16#0A#),
      688 => to_slv(opcode_type, 16#08#),
      689 => to_slv(opcode_type, 16#0B#),
      690 => to_slv(opcode_type, 16#0C#),
      691 => to_slv(opcode_type, 16#09#),
      692 => to_slv(opcode_type, 16#08#),
      693 => to_slv(opcode_type, 16#A3#),
      694 => to_slv(opcode_type, 16#E3#),
      695 => to_slv(opcode_type, 16#07#),
      696 => to_slv(opcode_type, 16#0D#),
      697 => to_slv(opcode_type, 16#0E#),
      698 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#08#),
      705 => to_slv(opcode_type, 16#09#),
      706 => to_slv(opcode_type, 16#06#),
      707 => to_slv(opcode_type, 16#08#),
      708 => to_slv(opcode_type, 16#0E#),
      709 => to_slv(opcode_type, 16#0F#),
      710 => to_slv(opcode_type, 16#02#),
      711 => to_slv(opcode_type, 16#0F#),
      712 => to_slv(opcode_type, 16#06#),
      713 => to_slv(opcode_type, 16#06#),
      714 => to_slv(opcode_type, 16#0A#),
      715 => to_slv(opcode_type, 16#0A#),
      716 => to_slv(opcode_type, 16#05#),
      717 => to_slv(opcode_type, 16#0C#),
      718 => to_slv(opcode_type, 16#07#),
      719 => to_slv(opcode_type, 16#06#),
      720 => to_slv(opcode_type, 16#02#),
      721 => to_slv(opcode_type, 16#0E#),
      722 => to_slv(opcode_type, 16#08#),
      723 => to_slv(opcode_type, 16#0C#),
      724 => to_slv(opcode_type, 16#0A#),
      725 => to_slv(opcode_type, 16#08#),
      726 => to_slv(opcode_type, 16#04#),
      727 => to_slv(opcode_type, 16#0B#),
      728 => to_slv(opcode_type, 16#04#),
      729 => to_slv(opcode_type, 16#10#),
      730 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#08#),
      737 => to_slv(opcode_type, 16#07#),
      738 => to_slv(opcode_type, 16#07#),
      739 => to_slv(opcode_type, 16#03#),
      740 => to_slv(opcode_type, 16#0A#),
      741 => to_slv(opcode_type, 16#07#),
      742 => to_slv(opcode_type, 16#0F#),
      743 => to_slv(opcode_type, 16#0B#),
      744 => to_slv(opcode_type, 16#01#),
      745 => to_slv(opcode_type, 16#03#),
      746 => to_slv(opcode_type, 16#11#),
      747 => to_slv(opcode_type, 16#07#),
      748 => to_slv(opcode_type, 16#07#),
      749 => to_slv(opcode_type, 16#09#),
      750 => to_slv(opcode_type, 16#39#),
      751 => to_slv(opcode_type, 16#0B#),
      752 => to_slv(opcode_type, 16#09#),
      753 => to_slv(opcode_type, 16#79#),
      754 => to_slv(opcode_type, 16#78#),
      755 => to_slv(opcode_type, 16#07#),
      756 => to_slv(opcode_type, 16#07#),
      757 => to_slv(opcode_type, 16#0C#),
      758 => to_slv(opcode_type, 16#0A#),
      759 => to_slv(opcode_type, 16#09#),
      760 => to_slv(opcode_type, 16#FC#),
      761 => to_slv(opcode_type, 16#0D#),
      762 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#09#),
      769 => to_slv(opcode_type, 16#07#),
      770 => to_slv(opcode_type, 16#07#),
      771 => to_slv(opcode_type, 16#02#),
      772 => to_slv(opcode_type, 16#0A#),
      773 => to_slv(opcode_type, 16#09#),
      774 => to_slv(opcode_type, 16#0C#),
      775 => to_slv(opcode_type, 16#0D#),
      776 => to_slv(opcode_type, 16#06#),
      777 => to_slv(opcode_type, 16#04#),
      778 => to_slv(opcode_type, 16#0A#),
      779 => to_slv(opcode_type, 16#02#),
      780 => to_slv(opcode_type, 16#0D#),
      781 => to_slv(opcode_type, 16#06#),
      782 => to_slv(opcode_type, 16#06#),
      783 => to_slv(opcode_type, 16#01#),
      784 => to_slv(opcode_type, 16#0F#),
      785 => to_slv(opcode_type, 16#07#),
      786 => to_slv(opcode_type, 16#0C#),
      787 => to_slv(opcode_type, 16#0F#),
      788 => to_slv(opcode_type, 16#06#),
      789 => to_slv(opcode_type, 16#08#),
      790 => to_slv(opcode_type, 16#0A#),
      791 => to_slv(opcode_type, 16#0F#),
      792 => to_slv(opcode_type, 16#02#),
      793 => to_slv(opcode_type, 16#11#),
      794 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#08#),
      801 => to_slv(opcode_type, 16#08#),
      802 => to_slv(opcode_type, 16#09#),
      803 => to_slv(opcode_type, 16#03#),
      804 => to_slv(opcode_type, 16#0A#),
      805 => to_slv(opcode_type, 16#02#),
      806 => to_slv(opcode_type, 16#2F#),
      807 => to_slv(opcode_type, 16#05#),
      808 => to_slv(opcode_type, 16#08#),
      809 => to_slv(opcode_type, 16#0B#),
      810 => to_slv(opcode_type, 16#FD#),
      811 => to_slv(opcode_type, 16#07#),
      812 => to_slv(opcode_type, 16#07#),
      813 => to_slv(opcode_type, 16#07#),
      814 => to_slv(opcode_type, 16#86#),
      815 => to_slv(opcode_type, 16#FF#),
      816 => to_slv(opcode_type, 16#09#),
      817 => to_slv(opcode_type, 16#0A#),
      818 => to_slv(opcode_type, 16#0D#),
      819 => to_slv(opcode_type, 16#06#),
      820 => to_slv(opcode_type, 16#07#),
      821 => to_slv(opcode_type, 16#10#),
      822 => to_slv(opcode_type, 16#11#),
      823 => to_slv(opcode_type, 16#06#),
      824 => to_slv(opcode_type, 16#0B#),
      825 => to_slv(opcode_type, 16#0B#),
      826 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#09#),
      833 => to_slv(opcode_type, 16#07#),
      834 => to_slv(opcode_type, 16#04#),
      835 => to_slv(opcode_type, 16#06#),
      836 => to_slv(opcode_type, 16#0F#),
      837 => to_slv(opcode_type, 16#11#),
      838 => to_slv(opcode_type, 16#08#),
      839 => to_slv(opcode_type, 16#08#),
      840 => to_slv(opcode_type, 16#D5#),
      841 => to_slv(opcode_type, 16#0C#),
      842 => to_slv(opcode_type, 16#01#),
      843 => to_slv(opcode_type, 16#0E#),
      844 => to_slv(opcode_type, 16#08#),
      845 => to_slv(opcode_type, 16#06#),
      846 => to_slv(opcode_type, 16#06#),
      847 => to_slv(opcode_type, 16#0A#),
      848 => to_slv(opcode_type, 16#0F#),
      849 => to_slv(opcode_type, 16#03#),
      850 => to_slv(opcode_type, 16#0E#),
      851 => to_slv(opcode_type, 16#09#),
      852 => to_slv(opcode_type, 16#08#),
      853 => to_slv(opcode_type, 16#0E#),
      854 => to_slv(opcode_type, 16#0E#),
      855 => to_slv(opcode_type, 16#06#),
      856 => to_slv(opcode_type, 16#0B#),
      857 => to_slv(opcode_type, 16#10#),
      858 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#06#),
      865 => to_slv(opcode_type, 16#07#),
      866 => to_slv(opcode_type, 16#08#),
      867 => to_slv(opcode_type, 16#08#),
      868 => to_slv(opcode_type, 16#11#),
      869 => to_slv(opcode_type, 16#11#),
      870 => to_slv(opcode_type, 16#07#),
      871 => to_slv(opcode_type, 16#0F#),
      872 => to_slv(opcode_type, 16#0F#),
      873 => to_slv(opcode_type, 16#01#),
      874 => to_slv(opcode_type, 16#07#),
      875 => to_slv(opcode_type, 16#0B#),
      876 => to_slv(opcode_type, 16#0B#),
      877 => to_slv(opcode_type, 16#07#),
      878 => to_slv(opcode_type, 16#08#),
      879 => to_slv(opcode_type, 16#02#),
      880 => to_slv(opcode_type, 16#0E#),
      881 => to_slv(opcode_type, 16#01#),
      882 => to_slv(opcode_type, 16#0C#),
      883 => to_slv(opcode_type, 16#08#),
      884 => to_slv(opcode_type, 16#07#),
      885 => to_slv(opcode_type, 16#37#),
      886 => to_slv(opcode_type, 16#11#),
      887 => to_slv(opcode_type, 16#08#),
      888 => to_slv(opcode_type, 16#0A#),
      889 => to_slv(opcode_type, 16#0A#),
      890 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#06#),
      898 => to_slv(opcode_type, 16#08#),
      899 => to_slv(opcode_type, 16#01#),
      900 => to_slv(opcode_type, 16#0D#),
      901 => to_slv(opcode_type, 16#04#),
      902 => to_slv(opcode_type, 16#0F#),
      903 => to_slv(opcode_type, 16#02#),
      904 => to_slv(opcode_type, 16#09#),
      905 => to_slv(opcode_type, 16#0B#),
      906 => to_slv(opcode_type, 16#0E#),
      907 => to_slv(opcode_type, 16#07#),
      908 => to_slv(opcode_type, 16#08#),
      909 => to_slv(opcode_type, 16#09#),
      910 => to_slv(opcode_type, 16#0E#),
      911 => to_slv(opcode_type, 16#10#),
      912 => to_slv(opcode_type, 16#06#),
      913 => to_slv(opcode_type, 16#0C#),
      914 => to_slv(opcode_type, 16#0C#),
      915 => to_slv(opcode_type, 16#08#),
      916 => to_slv(opcode_type, 16#06#),
      917 => to_slv(opcode_type, 16#0E#),
      918 => to_slv(opcode_type, 16#EB#),
      919 => to_slv(opcode_type, 16#09#),
      920 => to_slv(opcode_type, 16#0D#),
      921 => to_slv(opcode_type, 16#11#),
      922 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#09#),
      929 => to_slv(opcode_type, 16#08#),
      930 => to_slv(opcode_type, 16#07#),
      931 => to_slv(opcode_type, 16#05#),
      932 => to_slv(opcode_type, 16#0E#),
      933 => to_slv(opcode_type, 16#01#),
      934 => to_slv(opcode_type, 16#0E#),
      935 => to_slv(opcode_type, 16#06#),
      936 => to_slv(opcode_type, 16#02#),
      937 => to_slv(opcode_type, 16#0C#),
      938 => to_slv(opcode_type, 16#03#),
      939 => to_slv(opcode_type, 16#0C#),
      940 => to_slv(opcode_type, 16#06#),
      941 => to_slv(opcode_type, 16#09#),
      942 => to_slv(opcode_type, 16#06#),
      943 => to_slv(opcode_type, 16#0D#),
      944 => to_slv(opcode_type, 16#EA#),
      945 => to_slv(opcode_type, 16#05#),
      946 => to_slv(opcode_type, 16#7A#),
      947 => to_slv(opcode_type, 16#06#),
      948 => to_slv(opcode_type, 16#08#),
      949 => to_slv(opcode_type, 16#0F#),
      950 => to_slv(opcode_type, 16#0B#),
      951 => to_slv(opcode_type, 16#08#),
      952 => to_slv(opcode_type, 16#11#),
      953 => to_slv(opcode_type, 16#0B#),
      954 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#08#),
      962 => to_slv(opcode_type, 16#08#),
      963 => to_slv(opcode_type, 16#09#),
      964 => to_slv(opcode_type, 16#0B#),
      965 => to_slv(opcode_type, 16#11#),
      966 => to_slv(opcode_type, 16#09#),
      967 => to_slv(opcode_type, 16#10#),
      968 => to_slv(opcode_type, 16#0A#),
      969 => to_slv(opcode_type, 16#01#),
      970 => to_slv(opcode_type, 16#02#),
      971 => to_slv(opcode_type, 16#0E#),
      972 => to_slv(opcode_type, 16#08#),
      973 => to_slv(opcode_type, 16#06#),
      974 => to_slv(opcode_type, 16#07#),
      975 => to_slv(opcode_type, 16#0C#),
      976 => to_slv(opcode_type, 16#10#),
      977 => to_slv(opcode_type, 16#03#),
      978 => to_slv(opcode_type, 16#0E#),
      979 => to_slv(opcode_type, 16#06#),
      980 => to_slv(opcode_type, 16#06#),
      981 => to_slv(opcode_type, 16#10#),
      982 => to_slv(opcode_type, 16#0D#),
      983 => to_slv(opcode_type, 16#09#),
      984 => to_slv(opcode_type, 16#0F#),
      985 => to_slv(opcode_type, 16#0A#),
      986 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#06#),
      993 => to_slv(opcode_type, 16#06#),
      994 => to_slv(opcode_type, 16#08#),
      995 => to_slv(opcode_type, 16#09#),
      996 => to_slv(opcode_type, 16#0A#),
      997 => to_slv(opcode_type, 16#0B#),
      998 => to_slv(opcode_type, 16#06#),
      999 => to_slv(opcode_type, 16#81#),
      1000 => to_slv(opcode_type, 16#0E#),
      1001 => to_slv(opcode_type, 16#06#),
      1002 => to_slv(opcode_type, 16#07#),
      1003 => to_slv(opcode_type, 16#10#),
      1004 => to_slv(opcode_type, 16#0C#),
      1005 => to_slv(opcode_type, 16#03#),
      1006 => to_slv(opcode_type, 16#0B#),
      1007 => to_slv(opcode_type, 16#07#),
      1008 => to_slv(opcode_type, 16#08#),
      1009 => to_slv(opcode_type, 16#01#),
      1010 => to_slv(opcode_type, 16#0B#),
      1011 => to_slv(opcode_type, 16#08#),
      1012 => to_slv(opcode_type, 16#0A#),
      1013 => to_slv(opcode_type, 16#0F#),
      1014 => to_slv(opcode_type, 16#07#),
      1015 => to_slv(opcode_type, 16#04#),
      1016 => to_slv(opcode_type, 16#11#),
      1017 => to_slv(opcode_type, 16#11#),
      1018 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#09#),
      1025 => to_slv(opcode_type, 16#09#),
      1026 => to_slv(opcode_type, 16#05#),
      1027 => to_slv(opcode_type, 16#02#),
      1028 => to_slv(opcode_type, 16#0C#),
      1029 => to_slv(opcode_type, 16#06#),
      1030 => to_slv(opcode_type, 16#02#),
      1031 => to_slv(opcode_type, 16#11#),
      1032 => to_slv(opcode_type, 16#07#),
      1033 => to_slv(opcode_type, 16#0C#),
      1034 => to_slv(opcode_type, 16#0E#),
      1035 => to_slv(opcode_type, 16#09#),
      1036 => to_slv(opcode_type, 16#09#),
      1037 => to_slv(opcode_type, 16#07#),
      1038 => to_slv(opcode_type, 16#0E#),
      1039 => to_slv(opcode_type, 16#0E#),
      1040 => to_slv(opcode_type, 16#07#),
      1041 => to_slv(opcode_type, 16#EC#),
      1042 => to_slv(opcode_type, 16#0A#),
      1043 => to_slv(opcode_type, 16#06#),
      1044 => to_slv(opcode_type, 16#07#),
      1045 => to_slv(opcode_type, 16#10#),
      1046 => to_slv(opcode_type, 16#10#),
      1047 => to_slv(opcode_type, 16#08#),
      1048 => to_slv(opcode_type, 16#0E#),
      1049 => to_slv(opcode_type, 16#0F#),
      1050 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#09#),
      1057 => to_slv(opcode_type, 16#09#),
      1058 => to_slv(opcode_type, 16#02#),
      1059 => to_slv(opcode_type, 16#02#),
      1060 => to_slv(opcode_type, 16#0C#),
      1061 => to_slv(opcode_type, 16#07#),
      1062 => to_slv(opcode_type, 16#06#),
      1063 => to_slv(opcode_type, 16#0F#),
      1064 => to_slv(opcode_type, 16#C1#),
      1065 => to_slv(opcode_type, 16#06#),
      1066 => to_slv(opcode_type, 16#0F#),
      1067 => to_slv(opcode_type, 16#11#),
      1068 => to_slv(opcode_type, 16#08#),
      1069 => to_slv(opcode_type, 16#07#),
      1070 => to_slv(opcode_type, 16#02#),
      1071 => to_slv(opcode_type, 16#10#),
      1072 => to_slv(opcode_type, 16#09#),
      1073 => to_slv(opcode_type, 16#0F#),
      1074 => to_slv(opcode_type, 16#0E#),
      1075 => to_slv(opcode_type, 16#07#),
      1076 => to_slv(opcode_type, 16#06#),
      1077 => to_slv(opcode_type, 16#0F#),
      1078 => to_slv(opcode_type, 16#0C#),
      1079 => to_slv(opcode_type, 16#07#),
      1080 => to_slv(opcode_type, 16#10#),
      1081 => to_slv(opcode_type, 16#0A#),
      1082 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#09#),
      1089 => to_slv(opcode_type, 16#09#),
      1090 => to_slv(opcode_type, 16#05#),
      1091 => to_slv(opcode_type, 16#06#),
      1092 => to_slv(opcode_type, 16#0A#),
      1093 => to_slv(opcode_type, 16#11#),
      1094 => to_slv(opcode_type, 16#06#),
      1095 => to_slv(opcode_type, 16#06#),
      1096 => to_slv(opcode_type, 16#0C#),
      1097 => to_slv(opcode_type, 16#10#),
      1098 => to_slv(opcode_type, 16#04#),
      1099 => to_slv(opcode_type, 16#0A#),
      1100 => to_slv(opcode_type, 16#07#),
      1101 => to_slv(opcode_type, 16#07#),
      1102 => to_slv(opcode_type, 16#05#),
      1103 => to_slv(opcode_type, 16#42#),
      1104 => to_slv(opcode_type, 16#07#),
      1105 => to_slv(opcode_type, 16#52#),
      1106 => to_slv(opcode_type, 16#0E#),
      1107 => to_slv(opcode_type, 16#07#),
      1108 => to_slv(opcode_type, 16#08#),
      1109 => to_slv(opcode_type, 16#0B#),
      1110 => to_slv(opcode_type, 16#D4#),
      1111 => to_slv(opcode_type, 16#06#),
      1112 => to_slv(opcode_type, 16#0F#),
      1113 => to_slv(opcode_type, 16#0A#),
      1114 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#08#),
      1121 => to_slv(opcode_type, 16#06#),
      1122 => to_slv(opcode_type, 16#03#),
      1123 => to_slv(opcode_type, 16#09#),
      1124 => to_slv(opcode_type, 16#0A#),
      1125 => to_slv(opcode_type, 16#11#),
      1126 => to_slv(opcode_type, 16#08#),
      1127 => to_slv(opcode_type, 16#02#),
      1128 => to_slv(opcode_type, 16#0B#),
      1129 => to_slv(opcode_type, 16#05#),
      1130 => to_slv(opcode_type, 16#10#),
      1131 => to_slv(opcode_type, 16#08#),
      1132 => to_slv(opcode_type, 16#07#),
      1133 => to_slv(opcode_type, 16#06#),
      1134 => to_slv(opcode_type, 16#0D#),
      1135 => to_slv(opcode_type, 16#AE#),
      1136 => to_slv(opcode_type, 16#06#),
      1137 => to_slv(opcode_type, 16#0D#),
      1138 => to_slv(opcode_type, 16#0B#),
      1139 => to_slv(opcode_type, 16#08#),
      1140 => to_slv(opcode_type, 16#08#),
      1141 => to_slv(opcode_type, 16#0C#),
      1142 => to_slv(opcode_type, 16#11#),
      1143 => to_slv(opcode_type, 16#09#),
      1144 => to_slv(opcode_type, 16#0D#),
      1145 => to_slv(opcode_type, 16#84#),
      1146 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#06#),
      1153 => to_slv(opcode_type, 16#09#),
      1154 => to_slv(opcode_type, 16#01#),
      1155 => to_slv(opcode_type, 16#07#),
      1156 => to_slv(opcode_type, 16#11#),
      1157 => to_slv(opcode_type, 16#D3#),
      1158 => to_slv(opcode_type, 16#09#),
      1159 => to_slv(opcode_type, 16#02#),
      1160 => to_slv(opcode_type, 16#0F#),
      1161 => to_slv(opcode_type, 16#06#),
      1162 => to_slv(opcode_type, 16#78#),
      1163 => to_slv(opcode_type, 16#0E#),
      1164 => to_slv(opcode_type, 16#06#),
      1165 => to_slv(opcode_type, 16#06#),
      1166 => to_slv(opcode_type, 16#02#),
      1167 => to_slv(opcode_type, 16#DF#),
      1168 => to_slv(opcode_type, 16#07#),
      1169 => to_slv(opcode_type, 16#11#),
      1170 => to_slv(opcode_type, 16#11#),
      1171 => to_slv(opcode_type, 16#09#),
      1172 => to_slv(opcode_type, 16#07#),
      1173 => to_slv(opcode_type, 16#10#),
      1174 => to_slv(opcode_type, 16#11#),
      1175 => to_slv(opcode_type, 16#07#),
      1176 => to_slv(opcode_type, 16#C6#),
      1177 => to_slv(opcode_type, 16#26#),
      1178 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#07#),
      1185 => to_slv(opcode_type, 16#07#),
      1186 => to_slv(opcode_type, 16#04#),
      1187 => to_slv(opcode_type, 16#08#),
      1188 => to_slv(opcode_type, 16#10#),
      1189 => to_slv(opcode_type, 16#0B#),
      1190 => to_slv(opcode_type, 16#07#),
      1191 => to_slv(opcode_type, 16#04#),
      1192 => to_slv(opcode_type, 16#0C#),
      1193 => to_slv(opcode_type, 16#08#),
      1194 => to_slv(opcode_type, 16#0B#),
      1195 => to_slv(opcode_type, 16#0B#),
      1196 => to_slv(opcode_type, 16#07#),
      1197 => to_slv(opcode_type, 16#09#),
      1198 => to_slv(opcode_type, 16#03#),
      1199 => to_slv(opcode_type, 16#11#),
      1200 => to_slv(opcode_type, 16#09#),
      1201 => to_slv(opcode_type, 16#0C#),
      1202 => to_slv(opcode_type, 16#0F#),
      1203 => to_slv(opcode_type, 16#09#),
      1204 => to_slv(opcode_type, 16#06#),
      1205 => to_slv(opcode_type, 16#0D#),
      1206 => to_slv(opcode_type, 16#10#),
      1207 => to_slv(opcode_type, 16#08#),
      1208 => to_slv(opcode_type, 16#11#),
      1209 => to_slv(opcode_type, 16#72#),
      1210 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#08#),
      1217 => to_slv(opcode_type, 16#07#),
      1218 => to_slv(opcode_type, 16#09#),
      1219 => to_slv(opcode_type, 16#02#),
      1220 => to_slv(opcode_type, 16#0D#),
      1221 => to_slv(opcode_type, 16#07#),
      1222 => to_slv(opcode_type, 16#0F#),
      1223 => to_slv(opcode_type, 16#10#),
      1224 => to_slv(opcode_type, 16#04#),
      1225 => to_slv(opcode_type, 16#04#),
      1226 => to_slv(opcode_type, 16#10#),
      1227 => to_slv(opcode_type, 16#06#),
      1228 => to_slv(opcode_type, 16#08#),
      1229 => to_slv(opcode_type, 16#08#),
      1230 => to_slv(opcode_type, 16#0F#),
      1231 => to_slv(opcode_type, 16#0A#),
      1232 => to_slv(opcode_type, 16#07#),
      1233 => to_slv(opcode_type, 16#0B#),
      1234 => to_slv(opcode_type, 16#0D#),
      1235 => to_slv(opcode_type, 16#06#),
      1236 => to_slv(opcode_type, 16#07#),
      1237 => to_slv(opcode_type, 16#0E#),
      1238 => to_slv(opcode_type, 16#10#),
      1239 => to_slv(opcode_type, 16#07#),
      1240 => to_slv(opcode_type, 16#0D#),
      1241 => to_slv(opcode_type, 16#11#),
      1242 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#06#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#02#),
      1251 => to_slv(opcode_type, 16#09#),
      1252 => to_slv(opcode_type, 16#0D#),
      1253 => to_slv(opcode_type, 16#11#),
      1254 => to_slv(opcode_type, 16#06#),
      1255 => to_slv(opcode_type, 16#09#),
      1256 => to_slv(opcode_type, 16#0E#),
      1257 => to_slv(opcode_type, 16#0C#),
      1258 => to_slv(opcode_type, 16#01#),
      1259 => to_slv(opcode_type, 16#0C#),
      1260 => to_slv(opcode_type, 16#09#),
      1261 => to_slv(opcode_type, 16#07#),
      1262 => to_slv(opcode_type, 16#02#),
      1263 => to_slv(opcode_type, 16#0C#),
      1264 => to_slv(opcode_type, 16#07#),
      1265 => to_slv(opcode_type, 16#0B#),
      1266 => to_slv(opcode_type, 16#0E#),
      1267 => to_slv(opcode_type, 16#08#),
      1268 => to_slv(opcode_type, 16#09#),
      1269 => to_slv(opcode_type, 16#0D#),
      1270 => to_slv(opcode_type, 16#11#),
      1271 => to_slv(opcode_type, 16#09#),
      1272 => to_slv(opcode_type, 16#0D#),
      1273 => to_slv(opcode_type, 16#0F#),
      1274 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#06#),
      1281 => to_slv(opcode_type, 16#07#),
      1282 => to_slv(opcode_type, 16#06#),
      1283 => to_slv(opcode_type, 16#01#),
      1284 => to_slv(opcode_type, 16#79#),
      1285 => to_slv(opcode_type, 16#05#),
      1286 => to_slv(opcode_type, 16#0E#),
      1287 => to_slv(opcode_type, 16#01#),
      1288 => to_slv(opcode_type, 16#07#),
      1289 => to_slv(opcode_type, 16#10#),
      1290 => to_slv(opcode_type, 16#0A#),
      1291 => to_slv(opcode_type, 16#06#),
      1292 => to_slv(opcode_type, 16#08#),
      1293 => to_slv(opcode_type, 16#06#),
      1294 => to_slv(opcode_type, 16#0A#),
      1295 => to_slv(opcode_type, 16#0F#),
      1296 => to_slv(opcode_type, 16#09#),
      1297 => to_slv(opcode_type, 16#66#),
      1298 => to_slv(opcode_type, 16#0F#),
      1299 => to_slv(opcode_type, 16#06#),
      1300 => to_slv(opcode_type, 16#09#),
      1301 => to_slv(opcode_type, 16#0F#),
      1302 => to_slv(opcode_type, 16#0E#),
      1303 => to_slv(opcode_type, 16#09#),
      1304 => to_slv(opcode_type, 16#0A#),
      1305 => to_slv(opcode_type, 16#10#),
      1306 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#07#),
      1313 => to_slv(opcode_type, 16#09#),
      1314 => to_slv(opcode_type, 16#09#),
      1315 => to_slv(opcode_type, 16#01#),
      1316 => to_slv(opcode_type, 16#10#),
      1317 => to_slv(opcode_type, 16#08#),
      1318 => to_slv(opcode_type, 16#0B#),
      1319 => to_slv(opcode_type, 16#0D#),
      1320 => to_slv(opcode_type, 16#07#),
      1321 => to_slv(opcode_type, 16#01#),
      1322 => to_slv(opcode_type, 16#0D#),
      1323 => to_slv(opcode_type, 16#01#),
      1324 => to_slv(opcode_type, 16#0D#),
      1325 => to_slv(opcode_type, 16#06#),
      1326 => to_slv(opcode_type, 16#09#),
      1327 => to_slv(opcode_type, 16#06#),
      1328 => to_slv(opcode_type, 16#E2#),
      1329 => to_slv(opcode_type, 16#0B#),
      1330 => to_slv(opcode_type, 16#05#),
      1331 => to_slv(opcode_type, 16#11#),
      1332 => to_slv(opcode_type, 16#09#),
      1333 => to_slv(opcode_type, 16#08#),
      1334 => to_slv(opcode_type, 16#0C#),
      1335 => to_slv(opcode_type, 16#D3#),
      1336 => to_slv(opcode_type, 16#01#),
      1337 => to_slv(opcode_type, 16#0B#),
      1338 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#06#),
      1345 => to_slv(opcode_type, 16#09#),
      1346 => to_slv(opcode_type, 16#01#),
      1347 => to_slv(opcode_type, 16#07#),
      1348 => to_slv(opcode_type, 16#0E#),
      1349 => to_slv(opcode_type, 16#0D#),
      1350 => to_slv(opcode_type, 16#09#),
      1351 => to_slv(opcode_type, 16#01#),
      1352 => to_slv(opcode_type, 16#10#),
      1353 => to_slv(opcode_type, 16#07#),
      1354 => to_slv(opcode_type, 16#0E#),
      1355 => to_slv(opcode_type, 16#0C#),
      1356 => to_slv(opcode_type, 16#08#),
      1357 => to_slv(opcode_type, 16#09#),
      1358 => to_slv(opcode_type, 16#02#),
      1359 => to_slv(opcode_type, 16#0D#),
      1360 => to_slv(opcode_type, 16#07#),
      1361 => to_slv(opcode_type, 16#0C#),
      1362 => to_slv(opcode_type, 16#0B#),
      1363 => to_slv(opcode_type, 16#08#),
      1364 => to_slv(opcode_type, 16#07#),
      1365 => to_slv(opcode_type, 16#10#),
      1366 => to_slv(opcode_type, 16#0E#),
      1367 => to_slv(opcode_type, 16#08#),
      1368 => to_slv(opcode_type, 16#0C#),
      1369 => to_slv(opcode_type, 16#0F#),
      1370 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#06#),
      1377 => to_slv(opcode_type, 16#09#),
      1378 => to_slv(opcode_type, 16#09#),
      1379 => to_slv(opcode_type, 16#05#),
      1380 => to_slv(opcode_type, 16#10#),
      1381 => to_slv(opcode_type, 16#01#),
      1382 => to_slv(opcode_type, 16#11#),
      1383 => to_slv(opcode_type, 16#05#),
      1384 => to_slv(opcode_type, 16#07#),
      1385 => to_slv(opcode_type, 16#0D#),
      1386 => to_slv(opcode_type, 16#10#),
      1387 => to_slv(opcode_type, 16#07#),
      1388 => to_slv(opcode_type, 16#07#),
      1389 => to_slv(opcode_type, 16#08#),
      1390 => to_slv(opcode_type, 16#0C#),
      1391 => to_slv(opcode_type, 16#0A#),
      1392 => to_slv(opcode_type, 16#06#),
      1393 => to_slv(opcode_type, 16#41#),
      1394 => to_slv(opcode_type, 16#52#),
      1395 => to_slv(opcode_type, 16#06#),
      1396 => to_slv(opcode_type, 16#09#),
      1397 => to_slv(opcode_type, 16#10#),
      1398 => to_slv(opcode_type, 16#0E#),
      1399 => to_slv(opcode_type, 16#06#),
      1400 => to_slv(opcode_type, 16#0C#),
      1401 => to_slv(opcode_type, 16#11#),
      1402 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#09#),
      1410 => to_slv(opcode_type, 16#05#),
      1411 => to_slv(opcode_type, 16#02#),
      1412 => to_slv(opcode_type, 16#0C#),
      1413 => to_slv(opcode_type, 16#08#),
      1414 => to_slv(opcode_type, 16#08#),
      1415 => to_slv(opcode_type, 16#0F#),
      1416 => to_slv(opcode_type, 16#0A#),
      1417 => to_slv(opcode_type, 16#05#),
      1418 => to_slv(opcode_type, 16#0D#),
      1419 => to_slv(opcode_type, 16#07#),
      1420 => to_slv(opcode_type, 16#08#),
      1421 => to_slv(opcode_type, 16#06#),
      1422 => to_slv(opcode_type, 16#0E#),
      1423 => to_slv(opcode_type, 16#0B#),
      1424 => to_slv(opcode_type, 16#06#),
      1425 => to_slv(opcode_type, 16#0D#),
      1426 => to_slv(opcode_type, 16#0F#),
      1427 => to_slv(opcode_type, 16#08#),
      1428 => to_slv(opcode_type, 16#08#),
      1429 => to_slv(opcode_type, 16#0E#),
      1430 => to_slv(opcode_type, 16#0E#),
      1431 => to_slv(opcode_type, 16#07#),
      1432 => to_slv(opcode_type, 16#0B#),
      1433 => to_slv(opcode_type, 16#24#),
      1434 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#07#),
      1441 => to_slv(opcode_type, 16#07#),
      1442 => to_slv(opcode_type, 16#05#),
      1443 => to_slv(opcode_type, 16#02#),
      1444 => to_slv(opcode_type, 16#0A#),
      1445 => to_slv(opcode_type, 16#06#),
      1446 => to_slv(opcode_type, 16#02#),
      1447 => to_slv(opcode_type, 16#0C#),
      1448 => to_slv(opcode_type, 16#06#),
      1449 => to_slv(opcode_type, 16#11#),
      1450 => to_slv(opcode_type, 16#11#),
      1451 => to_slv(opcode_type, 16#06#),
      1452 => to_slv(opcode_type, 16#09#),
      1453 => to_slv(opcode_type, 16#07#),
      1454 => to_slv(opcode_type, 16#0B#),
      1455 => to_slv(opcode_type, 16#0D#),
      1456 => to_slv(opcode_type, 16#06#),
      1457 => to_slv(opcode_type, 16#88#),
      1458 => to_slv(opcode_type, 16#0D#),
      1459 => to_slv(opcode_type, 16#06#),
      1460 => to_slv(opcode_type, 16#08#),
      1461 => to_slv(opcode_type, 16#0B#),
      1462 => to_slv(opcode_type, 16#0D#),
      1463 => to_slv(opcode_type, 16#08#),
      1464 => to_slv(opcode_type, 16#0A#),
      1465 => to_slv(opcode_type, 16#0D#),
      1466 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#07#),
      1473 => to_slv(opcode_type, 16#07#),
      1474 => to_slv(opcode_type, 16#07#),
      1475 => to_slv(opcode_type, 16#05#),
      1476 => to_slv(opcode_type, 16#0F#),
      1477 => to_slv(opcode_type, 16#04#),
      1478 => to_slv(opcode_type, 16#0B#),
      1479 => to_slv(opcode_type, 16#08#),
      1480 => to_slv(opcode_type, 16#05#),
      1481 => to_slv(opcode_type, 16#0E#),
      1482 => to_slv(opcode_type, 16#05#),
      1483 => to_slv(opcode_type, 16#0C#),
      1484 => to_slv(opcode_type, 16#08#),
      1485 => to_slv(opcode_type, 16#07#),
      1486 => to_slv(opcode_type, 16#04#),
      1487 => to_slv(opcode_type, 16#6F#),
      1488 => to_slv(opcode_type, 16#06#),
      1489 => to_slv(opcode_type, 16#10#),
      1490 => to_slv(opcode_type, 16#0E#),
      1491 => to_slv(opcode_type, 16#07#),
      1492 => to_slv(opcode_type, 16#09#),
      1493 => to_slv(opcode_type, 16#0F#),
      1494 => to_slv(opcode_type, 16#10#),
      1495 => to_slv(opcode_type, 16#09#),
      1496 => to_slv(opcode_type, 16#0B#),
      1497 => to_slv(opcode_type, 16#0B#),
      1498 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#06#),
      1505 => to_slv(opcode_type, 16#08#),
      1506 => to_slv(opcode_type, 16#09#),
      1507 => to_slv(opcode_type, 16#06#),
      1508 => to_slv(opcode_type, 16#0D#),
      1509 => to_slv(opcode_type, 16#0B#),
      1510 => to_slv(opcode_type, 16#04#),
      1511 => to_slv(opcode_type, 16#0A#),
      1512 => to_slv(opcode_type, 16#02#),
      1513 => to_slv(opcode_type, 16#01#),
      1514 => to_slv(opcode_type, 16#0A#),
      1515 => to_slv(opcode_type, 16#08#),
      1516 => to_slv(opcode_type, 16#08#),
      1517 => to_slv(opcode_type, 16#07#),
      1518 => to_slv(opcode_type, 16#0F#),
      1519 => to_slv(opcode_type, 16#0E#),
      1520 => to_slv(opcode_type, 16#07#),
      1521 => to_slv(opcode_type, 16#11#),
      1522 => to_slv(opcode_type, 16#53#),
      1523 => to_slv(opcode_type, 16#07#),
      1524 => to_slv(opcode_type, 16#08#),
      1525 => to_slv(opcode_type, 16#11#),
      1526 => to_slv(opcode_type, 16#0E#),
      1527 => to_slv(opcode_type, 16#09#),
      1528 => to_slv(opcode_type, 16#10#),
      1529 => to_slv(opcode_type, 16#0D#),
      1530 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#06#),
      1537 => to_slv(opcode_type, 16#07#),
      1538 => to_slv(opcode_type, 16#06#),
      1539 => to_slv(opcode_type, 16#07#),
      1540 => to_slv(opcode_type, 16#10#),
      1541 => to_slv(opcode_type, 16#0D#),
      1542 => to_slv(opcode_type, 16#06#),
      1543 => to_slv(opcode_type, 16#0C#),
      1544 => to_slv(opcode_type, 16#11#),
      1545 => to_slv(opcode_type, 16#09#),
      1546 => to_slv(opcode_type, 16#04#),
      1547 => to_slv(opcode_type, 16#0D#),
      1548 => to_slv(opcode_type, 16#07#),
      1549 => to_slv(opcode_type, 16#0C#),
      1550 => to_slv(opcode_type, 16#10#),
      1551 => to_slv(opcode_type, 16#09#),
      1552 => to_slv(opcode_type, 16#08#),
      1553 => to_slv(opcode_type, 16#05#),
      1554 => to_slv(opcode_type, 16#0F#),
      1555 => to_slv(opcode_type, 16#08#),
      1556 => to_slv(opcode_type, 16#0D#),
      1557 => to_slv(opcode_type, 16#0C#),
      1558 => to_slv(opcode_type, 16#03#),
      1559 => to_slv(opcode_type, 16#07#),
      1560 => to_slv(opcode_type, 16#0F#),
      1561 => to_slv(opcode_type, 16#0D#),
      1562 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#09#),
      1569 => to_slv(opcode_type, 16#07#),
      1570 => to_slv(opcode_type, 16#07#),
      1571 => to_slv(opcode_type, 16#03#),
      1572 => to_slv(opcode_type, 16#0B#),
      1573 => to_slv(opcode_type, 16#04#),
      1574 => to_slv(opcode_type, 16#CB#),
      1575 => to_slv(opcode_type, 16#01#),
      1576 => to_slv(opcode_type, 16#08#),
      1577 => to_slv(opcode_type, 16#0D#),
      1578 => to_slv(opcode_type, 16#E9#),
      1579 => to_slv(opcode_type, 16#08#),
      1580 => to_slv(opcode_type, 16#07#),
      1581 => to_slv(opcode_type, 16#08#),
      1582 => to_slv(opcode_type, 16#11#),
      1583 => to_slv(opcode_type, 16#10#),
      1584 => to_slv(opcode_type, 16#07#),
      1585 => to_slv(opcode_type, 16#B4#),
      1586 => to_slv(opcode_type, 16#0A#),
      1587 => to_slv(opcode_type, 16#06#),
      1588 => to_slv(opcode_type, 16#08#),
      1589 => to_slv(opcode_type, 16#0D#),
      1590 => to_slv(opcode_type, 16#11#),
      1591 => to_slv(opcode_type, 16#09#),
      1592 => to_slv(opcode_type, 16#0F#),
      1593 => to_slv(opcode_type, 16#0C#),
      1594 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#07#),
      1602 => to_slv(opcode_type, 16#06#),
      1603 => to_slv(opcode_type, 16#08#),
      1604 => to_slv(opcode_type, 16#95#),
      1605 => to_slv(opcode_type, 16#0C#),
      1606 => to_slv(opcode_type, 16#07#),
      1607 => to_slv(opcode_type, 16#0B#),
      1608 => to_slv(opcode_type, 16#0C#),
      1609 => to_slv(opcode_type, 16#02#),
      1610 => to_slv(opcode_type, 16#02#),
      1611 => to_slv(opcode_type, 16#0F#),
      1612 => to_slv(opcode_type, 16#08#),
      1613 => to_slv(opcode_type, 16#09#),
      1614 => to_slv(opcode_type, 16#02#),
      1615 => to_slv(opcode_type, 16#10#),
      1616 => to_slv(opcode_type, 16#07#),
      1617 => to_slv(opcode_type, 16#0B#),
      1618 => to_slv(opcode_type, 16#0A#),
      1619 => to_slv(opcode_type, 16#08#),
      1620 => to_slv(opcode_type, 16#06#),
      1621 => to_slv(opcode_type, 16#0B#),
      1622 => to_slv(opcode_type, 16#0A#),
      1623 => to_slv(opcode_type, 16#08#),
      1624 => to_slv(opcode_type, 16#11#),
      1625 => to_slv(opcode_type, 16#99#),
      1626 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#07#),
      1633 => to_slv(opcode_type, 16#09#),
      1634 => to_slv(opcode_type, 16#07#),
      1635 => to_slv(opcode_type, 16#01#),
      1636 => to_slv(opcode_type, 16#0C#),
      1637 => to_slv(opcode_type, 16#02#),
      1638 => to_slv(opcode_type, 16#0D#),
      1639 => to_slv(opcode_type, 16#07#),
      1640 => to_slv(opcode_type, 16#01#),
      1641 => to_slv(opcode_type, 16#8D#),
      1642 => to_slv(opcode_type, 16#07#),
      1643 => to_slv(opcode_type, 16#0E#),
      1644 => to_slv(opcode_type, 16#0D#),
      1645 => to_slv(opcode_type, 16#07#),
      1646 => to_slv(opcode_type, 16#06#),
      1647 => to_slv(opcode_type, 16#06#),
      1648 => to_slv(opcode_type, 16#10#),
      1649 => to_slv(opcode_type, 16#BB#),
      1650 => to_slv(opcode_type, 16#03#),
      1651 => to_slv(opcode_type, 16#0C#),
      1652 => to_slv(opcode_type, 16#09#),
      1653 => to_slv(opcode_type, 16#06#),
      1654 => to_slv(opcode_type, 16#0E#),
      1655 => to_slv(opcode_type, 16#0A#),
      1656 => to_slv(opcode_type, 16#02#),
      1657 => to_slv(opcode_type, 16#0E#),
      1658 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#08#),
      1665 => to_slv(opcode_type, 16#08#),
      1666 => to_slv(opcode_type, 16#06#),
      1667 => to_slv(opcode_type, 16#03#),
      1668 => to_slv(opcode_type, 16#58#),
      1669 => to_slv(opcode_type, 16#04#),
      1670 => to_slv(opcode_type, 16#11#),
      1671 => to_slv(opcode_type, 16#02#),
      1672 => to_slv(opcode_type, 16#09#),
      1673 => to_slv(opcode_type, 16#0C#),
      1674 => to_slv(opcode_type, 16#11#),
      1675 => to_slv(opcode_type, 16#06#),
      1676 => to_slv(opcode_type, 16#09#),
      1677 => to_slv(opcode_type, 16#08#),
      1678 => to_slv(opcode_type, 16#10#),
      1679 => to_slv(opcode_type, 16#0D#),
      1680 => to_slv(opcode_type, 16#07#),
      1681 => to_slv(opcode_type, 16#0F#),
      1682 => to_slv(opcode_type, 16#0D#),
      1683 => to_slv(opcode_type, 16#09#),
      1684 => to_slv(opcode_type, 16#08#),
      1685 => to_slv(opcode_type, 16#B2#),
      1686 => to_slv(opcode_type, 16#11#),
      1687 => to_slv(opcode_type, 16#09#),
      1688 => to_slv(opcode_type, 16#0A#),
      1689 => to_slv(opcode_type, 16#0F#),
      1690 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#08#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#07#),
      1699 => to_slv(opcode_type, 16#06#),
      1700 => to_slv(opcode_type, 16#0C#),
      1701 => to_slv(opcode_type, 16#10#),
      1702 => to_slv(opcode_type, 16#05#),
      1703 => to_slv(opcode_type, 16#0F#),
      1704 => to_slv(opcode_type, 16#05#),
      1705 => to_slv(opcode_type, 16#06#),
      1706 => to_slv(opcode_type, 16#0A#),
      1707 => to_slv(opcode_type, 16#0A#),
      1708 => to_slv(opcode_type, 16#07#),
      1709 => to_slv(opcode_type, 16#06#),
      1710 => to_slv(opcode_type, 16#03#),
      1711 => to_slv(opcode_type, 16#D0#),
      1712 => to_slv(opcode_type, 16#08#),
      1713 => to_slv(opcode_type, 16#0C#),
      1714 => to_slv(opcode_type, 16#11#),
      1715 => to_slv(opcode_type, 16#07#),
      1716 => to_slv(opcode_type, 16#06#),
      1717 => to_slv(opcode_type, 16#0C#),
      1718 => to_slv(opcode_type, 16#0B#),
      1719 => to_slv(opcode_type, 16#09#),
      1720 => to_slv(opcode_type, 16#0A#),
      1721 => to_slv(opcode_type, 16#10#),
      1722 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#08#),
      1729 => to_slv(opcode_type, 16#08#),
      1730 => to_slv(opcode_type, 16#03#),
      1731 => to_slv(opcode_type, 16#04#),
      1732 => to_slv(opcode_type, 16#0A#),
      1733 => to_slv(opcode_type, 16#08#),
      1734 => to_slv(opcode_type, 16#04#),
      1735 => to_slv(opcode_type, 16#0E#),
      1736 => to_slv(opcode_type, 16#09#),
      1737 => to_slv(opcode_type, 16#11#),
      1738 => to_slv(opcode_type, 16#0E#),
      1739 => to_slv(opcode_type, 16#06#),
      1740 => to_slv(opcode_type, 16#06#),
      1741 => to_slv(opcode_type, 16#09#),
      1742 => to_slv(opcode_type, 16#0F#),
      1743 => to_slv(opcode_type, 16#10#),
      1744 => to_slv(opcode_type, 16#06#),
      1745 => to_slv(opcode_type, 16#11#),
      1746 => to_slv(opcode_type, 16#41#),
      1747 => to_slv(opcode_type, 16#07#),
      1748 => to_slv(opcode_type, 16#08#),
      1749 => to_slv(opcode_type, 16#0D#),
      1750 => to_slv(opcode_type, 16#10#),
      1751 => to_slv(opcode_type, 16#09#),
      1752 => to_slv(opcode_type, 16#0C#),
      1753 => to_slv(opcode_type, 16#0D#),
      1754 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#06#),
      1761 => to_slv(opcode_type, 16#09#),
      1762 => to_slv(opcode_type, 16#05#),
      1763 => to_slv(opcode_type, 16#06#),
      1764 => to_slv(opcode_type, 16#0F#),
      1765 => to_slv(opcode_type, 16#0C#),
      1766 => to_slv(opcode_type, 16#07#),
      1767 => to_slv(opcode_type, 16#09#),
      1768 => to_slv(opcode_type, 16#0E#),
      1769 => to_slv(opcode_type, 16#0E#),
      1770 => to_slv(opcode_type, 16#02#),
      1771 => to_slv(opcode_type, 16#85#),
      1772 => to_slv(opcode_type, 16#07#),
      1773 => to_slv(opcode_type, 16#06#),
      1774 => to_slv(opcode_type, 16#04#),
      1775 => to_slv(opcode_type, 16#58#),
      1776 => to_slv(opcode_type, 16#08#),
      1777 => to_slv(opcode_type, 16#BD#),
      1778 => to_slv(opcode_type, 16#0F#),
      1779 => to_slv(opcode_type, 16#09#),
      1780 => to_slv(opcode_type, 16#09#),
      1781 => to_slv(opcode_type, 16#10#),
      1782 => to_slv(opcode_type, 16#11#),
      1783 => to_slv(opcode_type, 16#09#),
      1784 => to_slv(opcode_type, 16#0F#),
      1785 => to_slv(opcode_type, 16#0F#),
      1786 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#06#),
      1793 => to_slv(opcode_type, 16#09#),
      1794 => to_slv(opcode_type, 16#06#),
      1795 => to_slv(opcode_type, 16#02#),
      1796 => to_slv(opcode_type, 16#11#),
      1797 => to_slv(opcode_type, 16#03#),
      1798 => to_slv(opcode_type, 16#10#),
      1799 => to_slv(opcode_type, 16#01#),
      1800 => to_slv(opcode_type, 16#08#),
      1801 => to_slv(opcode_type, 16#65#),
      1802 => to_slv(opcode_type, 16#0D#),
      1803 => to_slv(opcode_type, 16#07#),
      1804 => to_slv(opcode_type, 16#06#),
      1805 => to_slv(opcode_type, 16#09#),
      1806 => to_slv(opcode_type, 16#10#),
      1807 => to_slv(opcode_type, 16#10#),
      1808 => to_slv(opcode_type, 16#08#),
      1809 => to_slv(opcode_type, 16#11#),
      1810 => to_slv(opcode_type, 16#0A#),
      1811 => to_slv(opcode_type, 16#08#),
      1812 => to_slv(opcode_type, 16#07#),
      1813 => to_slv(opcode_type, 16#0F#),
      1814 => to_slv(opcode_type, 16#0C#),
      1815 => to_slv(opcode_type, 16#07#),
      1816 => to_slv(opcode_type, 16#0D#),
      1817 => to_slv(opcode_type, 16#0E#),
      1818 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#07#),
      1825 => to_slv(opcode_type, 16#08#),
      1826 => to_slv(opcode_type, 16#01#),
      1827 => to_slv(opcode_type, 16#08#),
      1828 => to_slv(opcode_type, 16#15#),
      1829 => to_slv(opcode_type, 16#0C#),
      1830 => to_slv(opcode_type, 16#06#),
      1831 => to_slv(opcode_type, 16#04#),
      1832 => to_slv(opcode_type, 16#0E#),
      1833 => to_slv(opcode_type, 16#01#),
      1834 => to_slv(opcode_type, 16#0A#),
      1835 => to_slv(opcode_type, 16#08#),
      1836 => to_slv(opcode_type, 16#07#),
      1837 => to_slv(opcode_type, 16#06#),
      1838 => to_slv(opcode_type, 16#10#),
      1839 => to_slv(opcode_type, 16#0B#),
      1840 => to_slv(opcode_type, 16#06#),
      1841 => to_slv(opcode_type, 16#0C#),
      1842 => to_slv(opcode_type, 16#0C#),
      1843 => to_slv(opcode_type, 16#06#),
      1844 => to_slv(opcode_type, 16#08#),
      1845 => to_slv(opcode_type, 16#0F#),
      1846 => to_slv(opcode_type, 16#10#),
      1847 => to_slv(opcode_type, 16#08#),
      1848 => to_slv(opcode_type, 16#0D#),
      1849 => to_slv(opcode_type, 16#0C#),
      1850 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#06#),
      1857 => to_slv(opcode_type, 16#09#),
      1858 => to_slv(opcode_type, 16#04#),
      1859 => to_slv(opcode_type, 16#05#),
      1860 => to_slv(opcode_type, 16#0D#),
      1861 => to_slv(opcode_type, 16#06#),
      1862 => to_slv(opcode_type, 16#09#),
      1863 => to_slv(opcode_type, 16#0C#),
      1864 => to_slv(opcode_type, 16#30#),
      1865 => to_slv(opcode_type, 16#01#),
      1866 => to_slv(opcode_type, 16#0C#),
      1867 => to_slv(opcode_type, 16#08#),
      1868 => to_slv(opcode_type, 16#06#),
      1869 => to_slv(opcode_type, 16#08#),
      1870 => to_slv(opcode_type, 16#0E#),
      1871 => to_slv(opcode_type, 16#11#),
      1872 => to_slv(opcode_type, 16#07#),
      1873 => to_slv(opcode_type, 16#0D#),
      1874 => to_slv(opcode_type, 16#7B#),
      1875 => to_slv(opcode_type, 16#06#),
      1876 => to_slv(opcode_type, 16#09#),
      1877 => to_slv(opcode_type, 16#0E#),
      1878 => to_slv(opcode_type, 16#0A#),
      1879 => to_slv(opcode_type, 16#06#),
      1880 => to_slv(opcode_type, 16#11#),
      1881 => to_slv(opcode_type, 16#11#),
      1882 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#08#),
      1890 => to_slv(opcode_type, 16#05#),
      1891 => to_slv(opcode_type, 16#06#),
      1892 => to_slv(opcode_type, 16#8C#),
      1893 => to_slv(opcode_type, 16#8D#),
      1894 => to_slv(opcode_type, 16#06#),
      1895 => to_slv(opcode_type, 16#05#),
      1896 => to_slv(opcode_type, 16#0D#),
      1897 => to_slv(opcode_type, 16#06#),
      1898 => to_slv(opcode_type, 16#CA#),
      1899 => to_slv(opcode_type, 16#0E#),
      1900 => to_slv(opcode_type, 16#07#),
      1901 => to_slv(opcode_type, 16#09#),
      1902 => to_slv(opcode_type, 16#06#),
      1903 => to_slv(opcode_type, 16#11#),
      1904 => to_slv(opcode_type, 16#0D#),
      1905 => to_slv(opcode_type, 16#02#),
      1906 => to_slv(opcode_type, 16#0B#),
      1907 => to_slv(opcode_type, 16#06#),
      1908 => to_slv(opcode_type, 16#09#),
      1909 => to_slv(opcode_type, 16#3D#),
      1910 => to_slv(opcode_type, 16#11#),
      1911 => to_slv(opcode_type, 16#09#),
      1912 => to_slv(opcode_type, 16#0E#),
      1913 => to_slv(opcode_type, 16#0C#),
      1914 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#09#),
      1921 => to_slv(opcode_type, 16#07#),
      1922 => to_slv(opcode_type, 16#05#),
      1923 => to_slv(opcode_type, 16#01#),
      1924 => to_slv(opcode_type, 16#10#),
      1925 => to_slv(opcode_type, 16#07#),
      1926 => to_slv(opcode_type, 16#09#),
      1927 => to_slv(opcode_type, 16#0E#),
      1928 => to_slv(opcode_type, 16#10#),
      1929 => to_slv(opcode_type, 16#07#),
      1930 => to_slv(opcode_type, 16#11#),
      1931 => to_slv(opcode_type, 16#10#),
      1932 => to_slv(opcode_type, 16#09#),
      1933 => to_slv(opcode_type, 16#06#),
      1934 => to_slv(opcode_type, 16#05#),
      1935 => to_slv(opcode_type, 16#0F#),
      1936 => to_slv(opcode_type, 16#07#),
      1937 => to_slv(opcode_type, 16#0A#),
      1938 => to_slv(opcode_type, 16#0D#),
      1939 => to_slv(opcode_type, 16#09#),
      1940 => to_slv(opcode_type, 16#08#),
      1941 => to_slv(opcode_type, 16#0B#),
      1942 => to_slv(opcode_type, 16#0F#),
      1943 => to_slv(opcode_type, 16#08#),
      1944 => to_slv(opcode_type, 16#0F#),
      1945 => to_slv(opcode_type, 16#0C#),
      1946 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#09#),
      1953 => to_slv(opcode_type, 16#08#),
      1954 => to_slv(opcode_type, 16#01#),
      1955 => to_slv(opcode_type, 16#04#),
      1956 => to_slv(opcode_type, 16#0D#),
      1957 => to_slv(opcode_type, 16#08#),
      1958 => to_slv(opcode_type, 16#03#),
      1959 => to_slv(opcode_type, 16#D6#),
      1960 => to_slv(opcode_type, 16#06#),
      1961 => to_slv(opcode_type, 16#0A#),
      1962 => to_slv(opcode_type, 16#AE#),
      1963 => to_slv(opcode_type, 16#09#),
      1964 => to_slv(opcode_type, 16#08#),
      1965 => to_slv(opcode_type, 16#06#),
      1966 => to_slv(opcode_type, 16#0C#),
      1967 => to_slv(opcode_type, 16#0F#),
      1968 => to_slv(opcode_type, 16#08#),
      1969 => to_slv(opcode_type, 16#0F#),
      1970 => to_slv(opcode_type, 16#0C#),
      1971 => to_slv(opcode_type, 16#07#),
      1972 => to_slv(opcode_type, 16#07#),
      1973 => to_slv(opcode_type, 16#0C#),
      1974 => to_slv(opcode_type, 16#0C#),
      1975 => to_slv(opcode_type, 16#08#),
      1976 => to_slv(opcode_type, 16#0F#),
      1977 => to_slv(opcode_type, 16#10#),
      1978 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#09#),
      1985 => to_slv(opcode_type, 16#09#),
      1986 => to_slv(opcode_type, 16#07#),
      1987 => to_slv(opcode_type, 16#01#),
      1988 => to_slv(opcode_type, 16#0D#),
      1989 => to_slv(opcode_type, 16#08#),
      1990 => to_slv(opcode_type, 16#0C#),
      1991 => to_slv(opcode_type, 16#0A#),
      1992 => to_slv(opcode_type, 16#06#),
      1993 => to_slv(opcode_type, 16#08#),
      1994 => to_slv(opcode_type, 16#11#),
      1995 => to_slv(opcode_type, 16#D0#),
      1996 => to_slv(opcode_type, 16#03#),
      1997 => to_slv(opcode_type, 16#0A#),
      1998 => to_slv(opcode_type, 16#07#),
      1999 => to_slv(opcode_type, 16#02#),
      2000 => to_slv(opcode_type, 16#09#),
      2001 => to_slv(opcode_type, 16#0F#),
      2002 => to_slv(opcode_type, 16#0E#),
      2003 => to_slv(opcode_type, 16#08#),
      2004 => to_slv(opcode_type, 16#08#),
      2005 => to_slv(opcode_type, 16#0A#),
      2006 => to_slv(opcode_type, 16#10#),
      2007 => to_slv(opcode_type, 16#09#),
      2008 => to_slv(opcode_type, 16#0B#),
      2009 => to_slv(opcode_type, 16#0F#),
      2010 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#07#),
      2017 => to_slv(opcode_type, 16#08#),
      2018 => to_slv(opcode_type, 16#07#),
      2019 => to_slv(opcode_type, 16#07#),
      2020 => to_slv(opcode_type, 16#0E#),
      2021 => to_slv(opcode_type, 16#0D#),
      2022 => to_slv(opcode_type, 16#02#),
      2023 => to_slv(opcode_type, 16#B8#),
      2024 => to_slv(opcode_type, 16#06#),
      2025 => to_slv(opcode_type, 16#08#),
      2026 => to_slv(opcode_type, 16#0F#),
      2027 => to_slv(opcode_type, 16#0D#),
      2028 => to_slv(opcode_type, 16#02#),
      2029 => to_slv(opcode_type, 16#0D#),
      2030 => to_slv(opcode_type, 16#07#),
      2031 => to_slv(opcode_type, 16#07#),
      2032 => to_slv(opcode_type, 16#01#),
      2033 => to_slv(opcode_type, 16#0C#),
      2034 => to_slv(opcode_type, 16#06#),
      2035 => to_slv(opcode_type, 16#8B#),
      2036 => to_slv(opcode_type, 16#0C#),
      2037 => to_slv(opcode_type, 16#08#),
      2038 => to_slv(opcode_type, 16#08#),
      2039 => to_slv(opcode_type, 16#0D#),
      2040 => to_slv(opcode_type, 16#0F#),
      2041 => to_slv(opcode_type, 16#0D#),
      2042 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#08#),
      2049 => to_slv(opcode_type, 16#07#),
      2050 => to_slv(opcode_type, 16#07#),
      2051 => to_slv(opcode_type, 16#02#),
      2052 => to_slv(opcode_type, 16#11#),
      2053 => to_slv(opcode_type, 16#06#),
      2054 => to_slv(opcode_type, 16#0F#),
      2055 => to_slv(opcode_type, 16#0F#),
      2056 => to_slv(opcode_type, 16#03#),
      2057 => to_slv(opcode_type, 16#04#),
      2058 => to_slv(opcode_type, 16#0F#),
      2059 => to_slv(opcode_type, 16#08#),
      2060 => to_slv(opcode_type, 16#09#),
      2061 => to_slv(opcode_type, 16#06#),
      2062 => to_slv(opcode_type, 16#0A#),
      2063 => to_slv(opcode_type, 16#FC#),
      2064 => to_slv(opcode_type, 16#09#),
      2065 => to_slv(opcode_type, 16#0A#),
      2066 => to_slv(opcode_type, 16#0B#),
      2067 => to_slv(opcode_type, 16#09#),
      2068 => to_slv(opcode_type, 16#07#),
      2069 => to_slv(opcode_type, 16#0B#),
      2070 => to_slv(opcode_type, 16#0E#),
      2071 => to_slv(opcode_type, 16#06#),
      2072 => to_slv(opcode_type, 16#0C#),
      2073 => to_slv(opcode_type, 16#11#),
      2074 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#09#),
      2081 => to_slv(opcode_type, 16#09#),
      2082 => to_slv(opcode_type, 16#08#),
      2083 => to_slv(opcode_type, 16#03#),
      2084 => to_slv(opcode_type, 16#0D#),
      2085 => to_slv(opcode_type, 16#08#),
      2086 => to_slv(opcode_type, 16#11#),
      2087 => to_slv(opcode_type, 16#0B#),
      2088 => to_slv(opcode_type, 16#06#),
      2089 => to_slv(opcode_type, 16#06#),
      2090 => to_slv(opcode_type, 16#11#),
      2091 => to_slv(opcode_type, 16#0F#),
      2092 => to_slv(opcode_type, 16#02#),
      2093 => to_slv(opcode_type, 16#0F#),
      2094 => to_slv(opcode_type, 16#07#),
      2095 => to_slv(opcode_type, 16#05#),
      2096 => to_slv(opcode_type, 16#09#),
      2097 => to_slv(opcode_type, 16#11#),
      2098 => to_slv(opcode_type, 16#10#),
      2099 => to_slv(opcode_type, 16#09#),
      2100 => to_slv(opcode_type, 16#06#),
      2101 => to_slv(opcode_type, 16#10#),
      2102 => to_slv(opcode_type, 16#10#),
      2103 => to_slv(opcode_type, 16#08#),
      2104 => to_slv(opcode_type, 16#0D#),
      2105 => to_slv(opcode_type, 16#0A#),
      2106 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#07#),
      2113 => to_slv(opcode_type, 16#07#),
      2114 => to_slv(opcode_type, 16#09#),
      2115 => to_slv(opcode_type, 16#07#),
      2116 => to_slv(opcode_type, 16#0B#),
      2117 => to_slv(opcode_type, 16#0F#),
      2118 => to_slv(opcode_type, 16#06#),
      2119 => to_slv(opcode_type, 16#0A#),
      2120 => to_slv(opcode_type, 16#0C#),
      2121 => to_slv(opcode_type, 16#09#),
      2122 => to_slv(opcode_type, 16#09#),
      2123 => to_slv(opcode_type, 16#0E#),
      2124 => to_slv(opcode_type, 16#0D#),
      2125 => to_slv(opcode_type, 16#01#),
      2126 => to_slv(opcode_type, 16#0E#),
      2127 => to_slv(opcode_type, 16#06#),
      2128 => to_slv(opcode_type, 16#04#),
      2129 => to_slv(opcode_type, 16#01#),
      2130 => to_slv(opcode_type, 16#0F#),
      2131 => to_slv(opcode_type, 16#07#),
      2132 => to_slv(opcode_type, 16#06#),
      2133 => to_slv(opcode_type, 16#11#),
      2134 => to_slv(opcode_type, 16#0D#),
      2135 => to_slv(opcode_type, 16#09#),
      2136 => to_slv(opcode_type, 16#11#),
      2137 => to_slv(opcode_type, 16#0D#),
      2138 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#08#),
      2146 => to_slv(opcode_type, 16#01#),
      2147 => to_slv(opcode_type, 16#02#),
      2148 => to_slv(opcode_type, 16#0C#),
      2149 => to_slv(opcode_type, 16#09#),
      2150 => to_slv(opcode_type, 16#07#),
      2151 => to_slv(opcode_type, 16#0A#),
      2152 => to_slv(opcode_type, 16#0E#),
      2153 => to_slv(opcode_type, 16#09#),
      2154 => to_slv(opcode_type, 16#10#),
      2155 => to_slv(opcode_type, 16#0F#),
      2156 => to_slv(opcode_type, 16#06#),
      2157 => to_slv(opcode_type, 16#06#),
      2158 => to_slv(opcode_type, 16#09#),
      2159 => to_slv(opcode_type, 16#10#),
      2160 => to_slv(opcode_type, 16#0B#),
      2161 => to_slv(opcode_type, 16#07#),
      2162 => to_slv(opcode_type, 16#28#),
      2163 => to_slv(opcode_type, 16#0D#),
      2164 => to_slv(opcode_type, 16#09#),
      2165 => to_slv(opcode_type, 16#01#),
      2166 => to_slv(opcode_type, 16#0C#),
      2167 => to_slv(opcode_type, 16#07#),
      2168 => to_slv(opcode_type, 16#0A#),
      2169 => to_slv(opcode_type, 16#0C#),
      2170 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#07#),
      2177 => to_slv(opcode_type, 16#09#),
      2178 => to_slv(opcode_type, 16#04#),
      2179 => to_slv(opcode_type, 16#04#),
      2180 => to_slv(opcode_type, 16#0E#),
      2181 => to_slv(opcode_type, 16#07#),
      2182 => to_slv(opcode_type, 16#02#),
      2183 => to_slv(opcode_type, 16#11#),
      2184 => to_slv(opcode_type, 16#07#),
      2185 => to_slv(opcode_type, 16#0E#),
      2186 => to_slv(opcode_type, 16#0A#),
      2187 => to_slv(opcode_type, 16#07#),
      2188 => to_slv(opcode_type, 16#07#),
      2189 => to_slv(opcode_type, 16#09#),
      2190 => to_slv(opcode_type, 16#0C#),
      2191 => to_slv(opcode_type, 16#0D#),
      2192 => to_slv(opcode_type, 16#08#),
      2193 => to_slv(opcode_type, 16#0C#),
      2194 => to_slv(opcode_type, 16#0E#),
      2195 => to_slv(opcode_type, 16#06#),
      2196 => to_slv(opcode_type, 16#07#),
      2197 => to_slv(opcode_type, 16#11#),
      2198 => to_slv(opcode_type, 16#DE#),
      2199 => to_slv(opcode_type, 16#07#),
      2200 => to_slv(opcode_type, 16#0F#),
      2201 => to_slv(opcode_type, 16#0E#),
      2202 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#08#),
      2209 => to_slv(opcode_type, 16#09#),
      2210 => to_slv(opcode_type, 16#05#),
      2211 => to_slv(opcode_type, 16#07#),
      2212 => to_slv(opcode_type, 16#11#),
      2213 => to_slv(opcode_type, 16#0D#),
      2214 => to_slv(opcode_type, 16#09#),
      2215 => to_slv(opcode_type, 16#03#),
      2216 => to_slv(opcode_type, 16#0E#),
      2217 => to_slv(opcode_type, 16#01#),
      2218 => to_slv(opcode_type, 16#0C#),
      2219 => to_slv(opcode_type, 16#08#),
      2220 => to_slv(opcode_type, 16#08#),
      2221 => to_slv(opcode_type, 16#08#),
      2222 => to_slv(opcode_type, 16#11#),
      2223 => to_slv(opcode_type, 16#0A#),
      2224 => to_slv(opcode_type, 16#09#),
      2225 => to_slv(opcode_type, 16#0B#),
      2226 => to_slv(opcode_type, 16#0D#),
      2227 => to_slv(opcode_type, 16#08#),
      2228 => to_slv(opcode_type, 16#09#),
      2229 => to_slv(opcode_type, 16#11#),
      2230 => to_slv(opcode_type, 16#0E#),
      2231 => to_slv(opcode_type, 16#09#),
      2232 => to_slv(opcode_type, 16#0E#),
      2233 => to_slv(opcode_type, 16#0D#),
      2234 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#07#),
      2241 => to_slv(opcode_type, 16#07#),
      2242 => to_slv(opcode_type, 16#05#),
      2243 => to_slv(opcode_type, 16#06#),
      2244 => to_slv(opcode_type, 16#10#),
      2245 => to_slv(opcode_type, 16#37#),
      2246 => to_slv(opcode_type, 16#09#),
      2247 => to_slv(opcode_type, 16#04#),
      2248 => to_slv(opcode_type, 16#11#),
      2249 => to_slv(opcode_type, 16#09#),
      2250 => to_slv(opcode_type, 16#11#),
      2251 => to_slv(opcode_type, 16#10#),
      2252 => to_slv(opcode_type, 16#06#),
      2253 => to_slv(opcode_type, 16#06#),
      2254 => to_slv(opcode_type, 16#06#),
      2255 => to_slv(opcode_type, 16#0A#),
      2256 => to_slv(opcode_type, 16#0D#),
      2257 => to_slv(opcode_type, 16#04#),
      2258 => to_slv(opcode_type, 16#11#),
      2259 => to_slv(opcode_type, 16#08#),
      2260 => to_slv(opcode_type, 16#06#),
      2261 => to_slv(opcode_type, 16#0C#),
      2262 => to_slv(opcode_type, 16#0F#),
      2263 => to_slv(opcode_type, 16#09#),
      2264 => to_slv(opcode_type, 16#0B#),
      2265 => to_slv(opcode_type, 16#0A#),
      2266 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#07#),
      2273 => to_slv(opcode_type, 16#07#),
      2274 => to_slv(opcode_type, 16#05#),
      2275 => to_slv(opcode_type, 16#02#),
      2276 => to_slv(opcode_type, 16#0D#),
      2277 => to_slv(opcode_type, 16#06#),
      2278 => to_slv(opcode_type, 16#01#),
      2279 => to_slv(opcode_type, 16#0C#),
      2280 => to_slv(opcode_type, 16#09#),
      2281 => to_slv(opcode_type, 16#0C#),
      2282 => to_slv(opcode_type, 16#8A#),
      2283 => to_slv(opcode_type, 16#09#),
      2284 => to_slv(opcode_type, 16#09#),
      2285 => to_slv(opcode_type, 16#09#),
      2286 => to_slv(opcode_type, 16#10#),
      2287 => to_slv(opcode_type, 16#43#),
      2288 => to_slv(opcode_type, 16#08#),
      2289 => to_slv(opcode_type, 16#0B#),
      2290 => to_slv(opcode_type, 16#0B#),
      2291 => to_slv(opcode_type, 16#08#),
      2292 => to_slv(opcode_type, 16#09#),
      2293 => to_slv(opcode_type, 16#0E#),
      2294 => to_slv(opcode_type, 16#0E#),
      2295 => to_slv(opcode_type, 16#06#),
      2296 => to_slv(opcode_type, 16#E7#),
      2297 => to_slv(opcode_type, 16#0D#),
      2298 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#09#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#09#),
      2307 => to_slv(opcode_type, 16#05#),
      2308 => to_slv(opcode_type, 16#0B#),
      2309 => to_slv(opcode_type, 16#07#),
      2310 => to_slv(opcode_type, 16#18#),
      2311 => to_slv(opcode_type, 16#10#),
      2312 => to_slv(opcode_type, 16#09#),
      2313 => to_slv(opcode_type, 16#08#),
      2314 => to_slv(opcode_type, 16#32#),
      2315 => to_slv(opcode_type, 16#0E#),
      2316 => to_slv(opcode_type, 16#01#),
      2317 => to_slv(opcode_type, 16#0C#),
      2318 => to_slv(opcode_type, 16#09#),
      2319 => to_slv(opcode_type, 16#03#),
      2320 => to_slv(opcode_type, 16#09#),
      2321 => to_slv(opcode_type, 16#10#),
      2322 => to_slv(opcode_type, 16#10#),
      2323 => to_slv(opcode_type, 16#09#),
      2324 => to_slv(opcode_type, 16#07#),
      2325 => to_slv(opcode_type, 16#0E#),
      2326 => to_slv(opcode_type, 16#0C#),
      2327 => to_slv(opcode_type, 16#09#),
      2328 => to_slv(opcode_type, 16#0A#),
      2329 => to_slv(opcode_type, 16#0A#),
      2330 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#07#),
      2337 => to_slv(opcode_type, 16#06#),
      2338 => to_slv(opcode_type, 16#09#),
      2339 => to_slv(opcode_type, 16#05#),
      2340 => to_slv(opcode_type, 16#0F#),
      2341 => to_slv(opcode_type, 16#06#),
      2342 => to_slv(opcode_type, 16#0B#),
      2343 => to_slv(opcode_type, 16#0A#),
      2344 => to_slv(opcode_type, 16#09#),
      2345 => to_slv(opcode_type, 16#06#),
      2346 => to_slv(opcode_type, 16#0D#),
      2347 => to_slv(opcode_type, 16#0F#),
      2348 => to_slv(opcode_type, 16#09#),
      2349 => to_slv(opcode_type, 16#0B#),
      2350 => to_slv(opcode_type, 16#10#),
      2351 => to_slv(opcode_type, 16#07#),
      2352 => to_slv(opcode_type, 16#04#),
      2353 => to_slv(opcode_type, 16#03#),
      2354 => to_slv(opcode_type, 16#14#),
      2355 => to_slv(opcode_type, 16#06#),
      2356 => to_slv(opcode_type, 16#07#),
      2357 => to_slv(opcode_type, 16#11#),
      2358 => to_slv(opcode_type, 16#0A#),
      2359 => to_slv(opcode_type, 16#09#),
      2360 => to_slv(opcode_type, 16#0A#),
      2361 => to_slv(opcode_type, 16#47#),
      2362 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#07#),
      2369 => to_slv(opcode_type, 16#07#),
      2370 => to_slv(opcode_type, 16#03#),
      2371 => to_slv(opcode_type, 16#09#),
      2372 => to_slv(opcode_type, 16#10#),
      2373 => to_slv(opcode_type, 16#0A#),
      2374 => to_slv(opcode_type, 16#06#),
      2375 => to_slv(opcode_type, 16#09#),
      2376 => to_slv(opcode_type, 16#0A#),
      2377 => to_slv(opcode_type, 16#10#),
      2378 => to_slv(opcode_type, 16#04#),
      2379 => to_slv(opcode_type, 16#0C#),
      2380 => to_slv(opcode_type, 16#06#),
      2381 => to_slv(opcode_type, 16#09#),
      2382 => to_slv(opcode_type, 16#09#),
      2383 => to_slv(opcode_type, 16#0D#),
      2384 => to_slv(opcode_type, 16#0A#),
      2385 => to_slv(opcode_type, 16#02#),
      2386 => to_slv(opcode_type, 16#8B#),
      2387 => to_slv(opcode_type, 16#06#),
      2388 => to_slv(opcode_type, 16#09#),
      2389 => to_slv(opcode_type, 16#0B#),
      2390 => to_slv(opcode_type, 16#0D#),
      2391 => to_slv(opcode_type, 16#07#),
      2392 => to_slv(opcode_type, 16#0F#),
      2393 => to_slv(opcode_type, 16#0C#),
      2394 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#08#),
      2401 => to_slv(opcode_type, 16#07#),
      2402 => to_slv(opcode_type, 16#01#),
      2403 => to_slv(opcode_type, 16#07#),
      2404 => to_slv(opcode_type, 16#10#),
      2405 => to_slv(opcode_type, 16#0B#),
      2406 => to_slv(opcode_type, 16#07#),
      2407 => to_slv(opcode_type, 16#02#),
      2408 => to_slv(opcode_type, 16#0F#),
      2409 => to_slv(opcode_type, 16#06#),
      2410 => to_slv(opcode_type, 16#14#),
      2411 => to_slv(opcode_type, 16#0F#),
      2412 => to_slv(opcode_type, 16#09#),
      2413 => to_slv(opcode_type, 16#08#),
      2414 => to_slv(opcode_type, 16#08#),
      2415 => to_slv(opcode_type, 16#0B#),
      2416 => to_slv(opcode_type, 16#11#),
      2417 => to_slv(opcode_type, 16#03#),
      2418 => to_slv(opcode_type, 16#10#),
      2419 => to_slv(opcode_type, 16#09#),
      2420 => to_slv(opcode_type, 16#08#),
      2421 => to_slv(opcode_type, 16#79#),
      2422 => to_slv(opcode_type, 16#0A#),
      2423 => to_slv(opcode_type, 16#08#),
      2424 => to_slv(opcode_type, 16#0C#),
      2425 => to_slv(opcode_type, 16#0E#),
      2426 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#07#),
      2433 => to_slv(opcode_type, 16#08#),
      2434 => to_slv(opcode_type, 16#01#),
      2435 => to_slv(opcode_type, 16#05#),
      2436 => to_slv(opcode_type, 16#11#),
      2437 => to_slv(opcode_type, 16#09#),
      2438 => to_slv(opcode_type, 16#03#),
      2439 => to_slv(opcode_type, 16#10#),
      2440 => to_slv(opcode_type, 16#09#),
      2441 => to_slv(opcode_type, 16#F0#),
      2442 => to_slv(opcode_type, 16#0E#),
      2443 => to_slv(opcode_type, 16#06#),
      2444 => to_slv(opcode_type, 16#09#),
      2445 => to_slv(opcode_type, 16#06#),
      2446 => to_slv(opcode_type, 16#0E#),
      2447 => to_slv(opcode_type, 16#0A#),
      2448 => to_slv(opcode_type, 16#06#),
      2449 => to_slv(opcode_type, 16#0C#),
      2450 => to_slv(opcode_type, 16#0C#),
      2451 => to_slv(opcode_type, 16#08#),
      2452 => to_slv(opcode_type, 16#09#),
      2453 => to_slv(opcode_type, 16#0D#),
      2454 => to_slv(opcode_type, 16#0D#),
      2455 => to_slv(opcode_type, 16#07#),
      2456 => to_slv(opcode_type, 16#0D#),
      2457 => to_slv(opcode_type, 16#11#),
      2458 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#09#),
      2465 => to_slv(opcode_type, 16#07#),
      2466 => to_slv(opcode_type, 16#08#),
      2467 => to_slv(opcode_type, 16#02#),
      2468 => to_slv(opcode_type, 16#0E#),
      2469 => to_slv(opcode_type, 16#07#),
      2470 => to_slv(opcode_type, 16#0E#),
      2471 => to_slv(opcode_type, 16#10#),
      2472 => to_slv(opcode_type, 16#06#),
      2473 => to_slv(opcode_type, 16#02#),
      2474 => to_slv(opcode_type, 16#0D#),
      2475 => to_slv(opcode_type, 16#02#),
      2476 => to_slv(opcode_type, 16#0B#),
      2477 => to_slv(opcode_type, 16#07#),
      2478 => to_slv(opcode_type, 16#07#),
      2479 => to_slv(opcode_type, 16#03#),
      2480 => to_slv(opcode_type, 16#10#),
      2481 => to_slv(opcode_type, 16#07#),
      2482 => to_slv(opcode_type, 16#0A#),
      2483 => to_slv(opcode_type, 16#0B#),
      2484 => to_slv(opcode_type, 16#07#),
      2485 => to_slv(opcode_type, 16#07#),
      2486 => to_slv(opcode_type, 16#0C#),
      2487 => to_slv(opcode_type, 16#11#),
      2488 => to_slv(opcode_type, 16#03#),
      2489 => to_slv(opcode_type, 16#0F#),
      2490 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#08#),
      2497 => to_slv(opcode_type, 16#08#),
      2498 => to_slv(opcode_type, 16#04#),
      2499 => to_slv(opcode_type, 16#09#),
      2500 => to_slv(opcode_type, 16#EE#),
      2501 => to_slv(opcode_type, 16#0F#),
      2502 => to_slv(opcode_type, 16#07#),
      2503 => to_slv(opcode_type, 16#05#),
      2504 => to_slv(opcode_type, 16#D4#),
      2505 => to_slv(opcode_type, 16#02#),
      2506 => to_slv(opcode_type, 16#0B#),
      2507 => to_slv(opcode_type, 16#09#),
      2508 => to_slv(opcode_type, 16#08#),
      2509 => to_slv(opcode_type, 16#07#),
      2510 => to_slv(opcode_type, 16#4D#),
      2511 => to_slv(opcode_type, 16#0B#),
      2512 => to_slv(opcode_type, 16#09#),
      2513 => to_slv(opcode_type, 16#10#),
      2514 => to_slv(opcode_type, 16#0C#),
      2515 => to_slv(opcode_type, 16#08#),
      2516 => to_slv(opcode_type, 16#09#),
      2517 => to_slv(opcode_type, 16#0C#),
      2518 => to_slv(opcode_type, 16#0D#),
      2519 => to_slv(opcode_type, 16#09#),
      2520 => to_slv(opcode_type, 16#10#),
      2521 => to_slv(opcode_type, 16#0D#),
      2522 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#06#),
      2530 => to_slv(opcode_type, 16#05#),
      2531 => to_slv(opcode_type, 16#07#),
      2532 => to_slv(opcode_type, 16#0B#),
      2533 => to_slv(opcode_type, 16#9D#),
      2534 => to_slv(opcode_type, 16#08#),
      2535 => to_slv(opcode_type, 16#04#),
      2536 => to_slv(opcode_type, 16#0B#),
      2537 => to_slv(opcode_type, 16#06#),
      2538 => to_slv(opcode_type, 16#0C#),
      2539 => to_slv(opcode_type, 16#0B#),
      2540 => to_slv(opcode_type, 16#06#),
      2541 => to_slv(opcode_type, 16#09#),
      2542 => to_slv(opcode_type, 16#03#),
      2543 => to_slv(opcode_type, 16#0B#),
      2544 => to_slv(opcode_type, 16#06#),
      2545 => to_slv(opcode_type, 16#0B#),
      2546 => to_slv(opcode_type, 16#98#),
      2547 => to_slv(opcode_type, 16#08#),
      2548 => to_slv(opcode_type, 16#07#),
      2549 => to_slv(opcode_type, 16#A7#),
      2550 => to_slv(opcode_type, 16#0D#),
      2551 => to_slv(opcode_type, 16#09#),
      2552 => to_slv(opcode_type, 16#17#),
      2553 => to_slv(opcode_type, 16#0F#),
      2554 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#08#),
      2561 => to_slv(opcode_type, 16#08#),
      2562 => to_slv(opcode_type, 16#08#),
      2563 => to_slv(opcode_type, 16#08#),
      2564 => to_slv(opcode_type, 16#10#),
      2565 => to_slv(opcode_type, 16#0E#),
      2566 => to_slv(opcode_type, 16#03#),
      2567 => to_slv(opcode_type, 16#0D#),
      2568 => to_slv(opcode_type, 16#06#),
      2569 => to_slv(opcode_type, 16#02#),
      2570 => to_slv(opcode_type, 16#0B#),
      2571 => to_slv(opcode_type, 16#01#),
      2572 => to_slv(opcode_type, 16#11#),
      2573 => to_slv(opcode_type, 16#06#),
      2574 => to_slv(opcode_type, 16#09#),
      2575 => to_slv(opcode_type, 16#03#),
      2576 => to_slv(opcode_type, 16#0C#),
      2577 => to_slv(opcode_type, 16#07#),
      2578 => to_slv(opcode_type, 16#0D#),
      2579 => to_slv(opcode_type, 16#0E#),
      2580 => to_slv(opcode_type, 16#09#),
      2581 => to_slv(opcode_type, 16#08#),
      2582 => to_slv(opcode_type, 16#0C#),
      2583 => to_slv(opcode_type, 16#11#),
      2584 => to_slv(opcode_type, 16#05#),
      2585 => to_slv(opcode_type, 16#0D#),
      2586 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#08#),
      2593 => to_slv(opcode_type, 16#06#),
      2594 => to_slv(opcode_type, 16#09#),
      2595 => to_slv(opcode_type, 16#05#),
      2596 => to_slv(opcode_type, 16#BC#),
      2597 => to_slv(opcode_type, 16#04#),
      2598 => to_slv(opcode_type, 16#0F#),
      2599 => to_slv(opcode_type, 16#08#),
      2600 => to_slv(opcode_type, 16#05#),
      2601 => to_slv(opcode_type, 16#0D#),
      2602 => to_slv(opcode_type, 16#06#),
      2603 => to_slv(opcode_type, 16#0D#),
      2604 => to_slv(opcode_type, 16#0B#),
      2605 => to_slv(opcode_type, 16#09#),
      2606 => to_slv(opcode_type, 16#09#),
      2607 => to_slv(opcode_type, 16#01#),
      2608 => to_slv(opcode_type, 16#0C#),
      2609 => to_slv(opcode_type, 16#03#),
      2610 => to_slv(opcode_type, 16#11#),
      2611 => to_slv(opcode_type, 16#06#),
      2612 => to_slv(opcode_type, 16#07#),
      2613 => to_slv(opcode_type, 16#0F#),
      2614 => to_slv(opcode_type, 16#0A#),
      2615 => to_slv(opcode_type, 16#06#),
      2616 => to_slv(opcode_type, 16#0D#),
      2617 => to_slv(opcode_type, 16#0B#),
      2618 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#09#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#06#),
      2627 => to_slv(opcode_type, 16#04#),
      2628 => to_slv(opcode_type, 16#0D#),
      2629 => to_slv(opcode_type, 16#08#),
      2630 => to_slv(opcode_type, 16#0C#),
      2631 => to_slv(opcode_type, 16#11#),
      2632 => to_slv(opcode_type, 16#05#),
      2633 => to_slv(opcode_type, 16#06#),
      2634 => to_slv(opcode_type, 16#0C#),
      2635 => to_slv(opcode_type, 16#0D#),
      2636 => to_slv(opcode_type, 16#08#),
      2637 => to_slv(opcode_type, 16#07#),
      2638 => to_slv(opcode_type, 16#09#),
      2639 => to_slv(opcode_type, 16#0A#),
      2640 => to_slv(opcode_type, 16#0F#),
      2641 => to_slv(opcode_type, 16#04#),
      2642 => to_slv(opcode_type, 16#0A#),
      2643 => to_slv(opcode_type, 16#07#),
      2644 => to_slv(opcode_type, 16#09#),
      2645 => to_slv(opcode_type, 16#0C#),
      2646 => to_slv(opcode_type, 16#0E#),
      2647 => to_slv(opcode_type, 16#09#),
      2648 => to_slv(opcode_type, 16#70#),
      2649 => to_slv(opcode_type, 16#10#),
      2650 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#06#),
      2657 => to_slv(opcode_type, 16#09#),
      2658 => to_slv(opcode_type, 16#08#),
      2659 => to_slv(opcode_type, 16#01#),
      2660 => to_slv(opcode_type, 16#0D#),
      2661 => to_slv(opcode_type, 16#03#),
      2662 => to_slv(opcode_type, 16#0D#),
      2663 => to_slv(opcode_type, 16#06#),
      2664 => to_slv(opcode_type, 16#07#),
      2665 => to_slv(opcode_type, 16#0C#),
      2666 => to_slv(opcode_type, 16#0F#),
      2667 => to_slv(opcode_type, 16#07#),
      2668 => to_slv(opcode_type, 16#0C#),
      2669 => to_slv(opcode_type, 16#0F#),
      2670 => to_slv(opcode_type, 16#08#),
      2671 => to_slv(opcode_type, 16#01#),
      2672 => to_slv(opcode_type, 16#09#),
      2673 => to_slv(opcode_type, 16#0C#),
      2674 => to_slv(opcode_type, 16#8E#),
      2675 => to_slv(opcode_type, 16#09#),
      2676 => to_slv(opcode_type, 16#08#),
      2677 => to_slv(opcode_type, 16#0C#),
      2678 => to_slv(opcode_type, 16#10#),
      2679 => to_slv(opcode_type, 16#08#),
      2680 => to_slv(opcode_type, 16#0A#),
      2681 => to_slv(opcode_type, 16#10#),
      2682 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#06#),
      2689 => to_slv(opcode_type, 16#08#),
      2690 => to_slv(opcode_type, 16#06#),
      2691 => to_slv(opcode_type, 16#06#),
      2692 => to_slv(opcode_type, 16#10#),
      2693 => to_slv(opcode_type, 16#0F#),
      2694 => to_slv(opcode_type, 16#08#),
      2695 => to_slv(opcode_type, 16#0E#),
      2696 => to_slv(opcode_type, 16#0A#),
      2697 => to_slv(opcode_type, 16#06#),
      2698 => to_slv(opcode_type, 16#08#),
      2699 => to_slv(opcode_type, 16#0D#),
      2700 => to_slv(opcode_type, 16#0E#),
      2701 => to_slv(opcode_type, 16#07#),
      2702 => to_slv(opcode_type, 16#0E#),
      2703 => to_slv(opcode_type, 16#0C#),
      2704 => to_slv(opcode_type, 16#09#),
      2705 => to_slv(opcode_type, 16#05#),
      2706 => to_slv(opcode_type, 16#09#),
      2707 => to_slv(opcode_type, 16#10#),
      2708 => to_slv(opcode_type, 16#0B#),
      2709 => to_slv(opcode_type, 16#07#),
      2710 => to_slv(opcode_type, 16#02#),
      2711 => to_slv(opcode_type, 16#0E#),
      2712 => to_slv(opcode_type, 16#05#),
      2713 => to_slv(opcode_type, 16#0E#),
      2714 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#06#),
      2721 => to_slv(opcode_type, 16#09#),
      2722 => to_slv(opcode_type, 16#08#),
      2723 => to_slv(opcode_type, 16#03#),
      2724 => to_slv(opcode_type, 16#0F#),
      2725 => to_slv(opcode_type, 16#09#),
      2726 => to_slv(opcode_type, 16#0B#),
      2727 => to_slv(opcode_type, 16#0E#),
      2728 => to_slv(opcode_type, 16#04#),
      2729 => to_slv(opcode_type, 16#03#),
      2730 => to_slv(opcode_type, 16#0D#),
      2731 => to_slv(opcode_type, 16#06#),
      2732 => to_slv(opcode_type, 16#06#),
      2733 => to_slv(opcode_type, 16#07#),
      2734 => to_slv(opcode_type, 16#0D#),
      2735 => to_slv(opcode_type, 16#0A#),
      2736 => to_slv(opcode_type, 16#08#),
      2737 => to_slv(opcode_type, 16#0D#),
      2738 => to_slv(opcode_type, 16#0D#),
      2739 => to_slv(opcode_type, 16#06#),
      2740 => to_slv(opcode_type, 16#09#),
      2741 => to_slv(opcode_type, 16#10#),
      2742 => to_slv(opcode_type, 16#0D#),
      2743 => to_slv(opcode_type, 16#08#),
      2744 => to_slv(opcode_type, 16#11#),
      2745 => to_slv(opcode_type, 16#11#),
      2746 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#06#),
      2753 => to_slv(opcode_type, 16#08#),
      2754 => to_slv(opcode_type, 16#04#),
      2755 => to_slv(opcode_type, 16#03#),
      2756 => to_slv(opcode_type, 16#2B#),
      2757 => to_slv(opcode_type, 16#07#),
      2758 => to_slv(opcode_type, 16#08#),
      2759 => to_slv(opcode_type, 16#0D#),
      2760 => to_slv(opcode_type, 16#0B#),
      2761 => to_slv(opcode_type, 16#07#),
      2762 => to_slv(opcode_type, 16#0B#),
      2763 => to_slv(opcode_type, 16#1C#),
      2764 => to_slv(opcode_type, 16#09#),
      2765 => to_slv(opcode_type, 16#06#),
      2766 => to_slv(opcode_type, 16#02#),
      2767 => to_slv(opcode_type, 16#0A#),
      2768 => to_slv(opcode_type, 16#07#),
      2769 => to_slv(opcode_type, 16#0A#),
      2770 => to_slv(opcode_type, 16#D1#),
      2771 => to_slv(opcode_type, 16#09#),
      2772 => to_slv(opcode_type, 16#07#),
      2773 => to_slv(opcode_type, 16#0F#),
      2774 => to_slv(opcode_type, 16#10#),
      2775 => to_slv(opcode_type, 16#07#),
      2776 => to_slv(opcode_type, 16#65#),
      2777 => to_slv(opcode_type, 16#0E#),
      2778 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#08#),
      2785 => to_slv(opcode_type, 16#09#),
      2786 => to_slv(opcode_type, 16#05#),
      2787 => to_slv(opcode_type, 16#07#),
      2788 => to_slv(opcode_type, 16#0C#),
      2789 => to_slv(opcode_type, 16#0F#),
      2790 => to_slv(opcode_type, 16#07#),
      2791 => to_slv(opcode_type, 16#06#),
      2792 => to_slv(opcode_type, 16#0C#),
      2793 => to_slv(opcode_type, 16#0A#),
      2794 => to_slv(opcode_type, 16#08#),
      2795 => to_slv(opcode_type, 16#0A#),
      2796 => to_slv(opcode_type, 16#0F#),
      2797 => to_slv(opcode_type, 16#07#),
      2798 => to_slv(opcode_type, 16#09#),
      2799 => to_slv(opcode_type, 16#07#),
      2800 => to_slv(opcode_type, 16#0B#),
      2801 => to_slv(opcode_type, 16#0E#),
      2802 => to_slv(opcode_type, 16#08#),
      2803 => to_slv(opcode_type, 16#0D#),
      2804 => to_slv(opcode_type, 16#0E#),
      2805 => to_slv(opcode_type, 16#09#),
      2806 => to_slv(opcode_type, 16#06#),
      2807 => to_slv(opcode_type, 16#0F#),
      2808 => to_slv(opcode_type, 16#10#),
      2809 => to_slv(opcode_type, 16#10#),
      2810 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#06#),
      2817 => to_slv(opcode_type, 16#09#),
      2818 => to_slv(opcode_type, 16#07#),
      2819 => to_slv(opcode_type, 16#09#),
      2820 => to_slv(opcode_type, 16#0A#),
      2821 => to_slv(opcode_type, 16#0D#),
      2822 => to_slv(opcode_type, 16#05#),
      2823 => to_slv(opcode_type, 16#0E#),
      2824 => to_slv(opcode_type, 16#06#),
      2825 => to_slv(opcode_type, 16#04#),
      2826 => to_slv(opcode_type, 16#0E#),
      2827 => to_slv(opcode_type, 16#04#),
      2828 => to_slv(opcode_type, 16#0E#),
      2829 => to_slv(opcode_type, 16#07#),
      2830 => to_slv(opcode_type, 16#07#),
      2831 => to_slv(opcode_type, 16#07#),
      2832 => to_slv(opcode_type, 16#0A#),
      2833 => to_slv(opcode_type, 16#0F#),
      2834 => to_slv(opcode_type, 16#06#),
      2835 => to_slv(opcode_type, 16#0A#),
      2836 => to_slv(opcode_type, 16#0F#),
      2837 => to_slv(opcode_type, 16#09#),
      2838 => to_slv(opcode_type, 16#02#),
      2839 => to_slv(opcode_type, 16#22#),
      2840 => to_slv(opcode_type, 16#02#),
      2841 => to_slv(opcode_type, 16#0E#),
      2842 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#07#),
      2849 => to_slv(opcode_type, 16#07#),
      2850 => to_slv(opcode_type, 16#03#),
      2851 => to_slv(opcode_type, 16#09#),
      2852 => to_slv(opcode_type, 16#0D#),
      2853 => to_slv(opcode_type, 16#0F#),
      2854 => to_slv(opcode_type, 16#06#),
      2855 => to_slv(opcode_type, 16#04#),
      2856 => to_slv(opcode_type, 16#11#),
      2857 => to_slv(opcode_type, 16#02#),
      2858 => to_slv(opcode_type, 16#3A#),
      2859 => to_slv(opcode_type, 16#08#),
      2860 => to_slv(opcode_type, 16#09#),
      2861 => to_slv(opcode_type, 16#08#),
      2862 => to_slv(opcode_type, 16#10#),
      2863 => to_slv(opcode_type, 16#12#),
      2864 => to_slv(opcode_type, 16#08#),
      2865 => to_slv(opcode_type, 16#11#),
      2866 => to_slv(opcode_type, 16#10#),
      2867 => to_slv(opcode_type, 16#07#),
      2868 => to_slv(opcode_type, 16#08#),
      2869 => to_slv(opcode_type, 16#2F#),
      2870 => to_slv(opcode_type, 16#10#),
      2871 => to_slv(opcode_type, 16#09#),
      2872 => to_slv(opcode_type, 16#0D#),
      2873 => to_slv(opcode_type, 16#0E#),
      2874 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#09#),
      2881 => to_slv(opcode_type, 16#06#),
      2882 => to_slv(opcode_type, 16#02#),
      2883 => to_slv(opcode_type, 16#08#),
      2884 => to_slv(opcode_type, 16#10#),
      2885 => to_slv(opcode_type, 16#10#),
      2886 => to_slv(opcode_type, 16#07#),
      2887 => to_slv(opcode_type, 16#02#),
      2888 => to_slv(opcode_type, 16#0D#),
      2889 => to_slv(opcode_type, 16#09#),
      2890 => to_slv(opcode_type, 16#0F#),
      2891 => to_slv(opcode_type, 16#0B#),
      2892 => to_slv(opcode_type, 16#08#),
      2893 => to_slv(opcode_type, 16#07#),
      2894 => to_slv(opcode_type, 16#05#),
      2895 => to_slv(opcode_type, 16#B0#),
      2896 => to_slv(opcode_type, 16#06#),
      2897 => to_slv(opcode_type, 16#0E#),
      2898 => to_slv(opcode_type, 16#0C#),
      2899 => to_slv(opcode_type, 16#07#),
      2900 => to_slv(opcode_type, 16#09#),
      2901 => to_slv(opcode_type, 16#10#),
      2902 => to_slv(opcode_type, 16#0B#),
      2903 => to_slv(opcode_type, 16#06#),
      2904 => to_slv(opcode_type, 16#0B#),
      2905 => to_slv(opcode_type, 16#25#),
      2906 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#08#),
      2913 => to_slv(opcode_type, 16#06#),
      2914 => to_slv(opcode_type, 16#06#),
      2915 => to_slv(opcode_type, 16#06#),
      2916 => to_slv(opcode_type, 16#0A#),
      2917 => to_slv(opcode_type, 16#0E#),
      2918 => to_slv(opcode_type, 16#04#),
      2919 => to_slv(opcode_type, 16#10#),
      2920 => to_slv(opcode_type, 16#08#),
      2921 => to_slv(opcode_type, 16#01#),
      2922 => to_slv(opcode_type, 16#11#),
      2923 => to_slv(opcode_type, 16#05#),
      2924 => to_slv(opcode_type, 16#0B#),
      2925 => to_slv(opcode_type, 16#08#),
      2926 => to_slv(opcode_type, 16#08#),
      2927 => to_slv(opcode_type, 16#02#),
      2928 => to_slv(opcode_type, 16#0E#),
      2929 => to_slv(opcode_type, 16#04#),
      2930 => to_slv(opcode_type, 16#11#),
      2931 => to_slv(opcode_type, 16#07#),
      2932 => to_slv(opcode_type, 16#09#),
      2933 => to_slv(opcode_type, 16#0F#),
      2934 => to_slv(opcode_type, 16#F1#),
      2935 => to_slv(opcode_type, 16#06#),
      2936 => to_slv(opcode_type, 16#10#),
      2937 => to_slv(opcode_type, 16#B0#),
      2938 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#07#),
      2945 => to_slv(opcode_type, 16#06#),
      2946 => to_slv(opcode_type, 16#06#),
      2947 => to_slv(opcode_type, 16#02#),
      2948 => to_slv(opcode_type, 16#0B#),
      2949 => to_slv(opcode_type, 16#09#),
      2950 => to_slv(opcode_type, 16#11#),
      2951 => to_slv(opcode_type, 16#CE#),
      2952 => to_slv(opcode_type, 16#05#),
      2953 => to_slv(opcode_type, 16#07#),
      2954 => to_slv(opcode_type, 16#0A#),
      2955 => to_slv(opcode_type, 16#10#),
      2956 => to_slv(opcode_type, 16#07#),
      2957 => to_slv(opcode_type, 16#06#),
      2958 => to_slv(opcode_type, 16#06#),
      2959 => to_slv(opcode_type, 16#E6#),
      2960 => to_slv(opcode_type, 16#0B#),
      2961 => to_slv(opcode_type, 16#05#),
      2962 => to_slv(opcode_type, 16#B7#),
      2963 => to_slv(opcode_type, 16#07#),
      2964 => to_slv(opcode_type, 16#08#),
      2965 => to_slv(opcode_type, 16#11#),
      2966 => to_slv(opcode_type, 16#11#),
      2967 => to_slv(opcode_type, 16#06#),
      2968 => to_slv(opcode_type, 16#0F#),
      2969 => to_slv(opcode_type, 16#0E#),
      2970 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#07#),
      2977 => to_slv(opcode_type, 16#08#),
      2978 => to_slv(opcode_type, 16#04#),
      2979 => to_slv(opcode_type, 16#09#),
      2980 => to_slv(opcode_type, 16#0D#),
      2981 => to_slv(opcode_type, 16#5B#),
      2982 => to_slv(opcode_type, 16#09#),
      2983 => to_slv(opcode_type, 16#02#),
      2984 => to_slv(opcode_type, 16#11#),
      2985 => to_slv(opcode_type, 16#09#),
      2986 => to_slv(opcode_type, 16#0A#),
      2987 => to_slv(opcode_type, 16#0D#),
      2988 => to_slv(opcode_type, 16#06#),
      2989 => to_slv(opcode_type, 16#07#),
      2990 => to_slv(opcode_type, 16#08#),
      2991 => to_slv(opcode_type, 16#0F#),
      2992 => to_slv(opcode_type, 16#11#),
      2993 => to_slv(opcode_type, 16#05#),
      2994 => to_slv(opcode_type, 16#0C#),
      2995 => to_slv(opcode_type, 16#07#),
      2996 => to_slv(opcode_type, 16#07#),
      2997 => to_slv(opcode_type, 16#0C#),
      2998 => to_slv(opcode_type, 16#0E#),
      2999 => to_slv(opcode_type, 16#06#),
      3000 => to_slv(opcode_type, 16#11#),
      3001 => to_slv(opcode_type, 16#C0#),
      3002 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#09#),
      3009 => to_slv(opcode_type, 16#09#),
      3010 => to_slv(opcode_type, 16#05#),
      3011 => to_slv(opcode_type, 16#06#),
      3012 => to_slv(opcode_type, 16#0D#),
      3013 => to_slv(opcode_type, 16#A5#),
      3014 => to_slv(opcode_type, 16#08#),
      3015 => to_slv(opcode_type, 16#06#),
      3016 => to_slv(opcode_type, 16#AB#),
      3017 => to_slv(opcode_type, 16#11#),
      3018 => to_slv(opcode_type, 16#01#),
      3019 => to_slv(opcode_type, 16#11#),
      3020 => to_slv(opcode_type, 16#07#),
      3021 => to_slv(opcode_type, 16#07#),
      3022 => to_slv(opcode_type, 16#03#),
      3023 => to_slv(opcode_type, 16#0B#),
      3024 => to_slv(opcode_type, 16#06#),
      3025 => to_slv(opcode_type, 16#11#),
      3026 => to_slv(opcode_type, 16#0E#),
      3027 => to_slv(opcode_type, 16#08#),
      3028 => to_slv(opcode_type, 16#06#),
      3029 => to_slv(opcode_type, 16#0B#),
      3030 => to_slv(opcode_type, 16#10#),
      3031 => to_slv(opcode_type, 16#06#),
      3032 => to_slv(opcode_type, 16#0B#),
      3033 => to_slv(opcode_type, 16#0D#),
      3034 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#07#),
      3041 => to_slv(opcode_type, 16#06#),
      3042 => to_slv(opcode_type, 16#01#),
      3043 => to_slv(opcode_type, 16#02#),
      3044 => to_slv(opcode_type, 16#0E#),
      3045 => to_slv(opcode_type, 16#09#),
      3046 => to_slv(opcode_type, 16#01#),
      3047 => to_slv(opcode_type, 16#0C#),
      3048 => to_slv(opcode_type, 16#08#),
      3049 => to_slv(opcode_type, 16#0A#),
      3050 => to_slv(opcode_type, 16#0D#),
      3051 => to_slv(opcode_type, 16#06#),
      3052 => to_slv(opcode_type, 16#08#),
      3053 => to_slv(opcode_type, 16#06#),
      3054 => to_slv(opcode_type, 16#0E#),
      3055 => to_slv(opcode_type, 16#0D#),
      3056 => to_slv(opcode_type, 16#08#),
      3057 => to_slv(opcode_type, 16#0B#),
      3058 => to_slv(opcode_type, 16#0B#),
      3059 => to_slv(opcode_type, 16#07#),
      3060 => to_slv(opcode_type, 16#06#),
      3061 => to_slv(opcode_type, 16#26#),
      3062 => to_slv(opcode_type, 16#0A#),
      3063 => to_slv(opcode_type, 16#08#),
      3064 => to_slv(opcode_type, 16#0C#),
      3065 => to_slv(opcode_type, 16#0E#),
      3066 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#08#),
      3073 => to_slv(opcode_type, 16#07#),
      3074 => to_slv(opcode_type, 16#07#),
      3075 => to_slv(opcode_type, 16#05#),
      3076 => to_slv(opcode_type, 16#10#),
      3077 => to_slv(opcode_type, 16#04#),
      3078 => to_slv(opcode_type, 16#11#),
      3079 => to_slv(opcode_type, 16#01#),
      3080 => to_slv(opcode_type, 16#07#),
      3081 => to_slv(opcode_type, 16#0B#),
      3082 => to_slv(opcode_type, 16#11#),
      3083 => to_slv(opcode_type, 16#08#),
      3084 => to_slv(opcode_type, 16#08#),
      3085 => to_slv(opcode_type, 16#08#),
      3086 => to_slv(opcode_type, 16#0C#),
      3087 => to_slv(opcode_type, 16#0F#),
      3088 => to_slv(opcode_type, 16#09#),
      3089 => to_slv(opcode_type, 16#0E#),
      3090 => to_slv(opcode_type, 16#11#),
      3091 => to_slv(opcode_type, 16#06#),
      3092 => to_slv(opcode_type, 16#09#),
      3093 => to_slv(opcode_type, 16#10#),
      3094 => to_slv(opcode_type, 16#0C#),
      3095 => to_slv(opcode_type, 16#06#),
      3096 => to_slv(opcode_type, 16#11#),
      3097 => to_slv(opcode_type, 16#70#),
      3098 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#08#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#03#),
      3107 => to_slv(opcode_type, 16#03#),
      3108 => to_slv(opcode_type, 16#92#),
      3109 => to_slv(opcode_type, 16#06#),
      3110 => to_slv(opcode_type, 16#09#),
      3111 => to_slv(opcode_type, 16#0D#),
      3112 => to_slv(opcode_type, 16#0A#),
      3113 => to_slv(opcode_type, 16#08#),
      3114 => to_slv(opcode_type, 16#0E#),
      3115 => to_slv(opcode_type, 16#75#),
      3116 => to_slv(opcode_type, 16#07#),
      3117 => to_slv(opcode_type, 16#06#),
      3118 => to_slv(opcode_type, 16#02#),
      3119 => to_slv(opcode_type, 16#0F#),
      3120 => to_slv(opcode_type, 16#08#),
      3121 => to_slv(opcode_type, 16#0D#),
      3122 => to_slv(opcode_type, 16#0F#),
      3123 => to_slv(opcode_type, 16#06#),
      3124 => to_slv(opcode_type, 16#09#),
      3125 => to_slv(opcode_type, 16#10#),
      3126 => to_slv(opcode_type, 16#0C#),
      3127 => to_slv(opcode_type, 16#09#),
      3128 => to_slv(opcode_type, 16#0B#),
      3129 => to_slv(opcode_type, 16#0B#),
      3130 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#07#),
      3137 => to_slv(opcode_type, 16#07#),
      3138 => to_slv(opcode_type, 16#03#),
      3139 => to_slv(opcode_type, 16#03#),
      3140 => to_slv(opcode_type, 16#0E#),
      3141 => to_slv(opcode_type, 16#09#),
      3142 => to_slv(opcode_type, 16#02#),
      3143 => to_slv(opcode_type, 16#0D#),
      3144 => to_slv(opcode_type, 16#08#),
      3145 => to_slv(opcode_type, 16#0F#),
      3146 => to_slv(opcode_type, 16#0C#),
      3147 => to_slv(opcode_type, 16#06#),
      3148 => to_slv(opcode_type, 16#09#),
      3149 => to_slv(opcode_type, 16#06#),
      3150 => to_slv(opcode_type, 16#0D#),
      3151 => to_slv(opcode_type, 16#0B#),
      3152 => to_slv(opcode_type, 16#08#),
      3153 => to_slv(opcode_type, 16#6D#),
      3154 => to_slv(opcode_type, 16#0D#),
      3155 => to_slv(opcode_type, 16#06#),
      3156 => to_slv(opcode_type, 16#07#),
      3157 => to_slv(opcode_type, 16#0D#),
      3158 => to_slv(opcode_type, 16#0D#),
      3159 => to_slv(opcode_type, 16#09#),
      3160 => to_slv(opcode_type, 16#11#),
      3161 => to_slv(opcode_type, 16#0A#),
      3162 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#07#),
      3169 => to_slv(opcode_type, 16#09#),
      3170 => to_slv(opcode_type, 16#02#),
      3171 => to_slv(opcode_type, 16#08#),
      3172 => to_slv(opcode_type, 16#10#),
      3173 => to_slv(opcode_type, 16#0D#),
      3174 => to_slv(opcode_type, 16#06#),
      3175 => to_slv(opcode_type, 16#08#),
      3176 => to_slv(opcode_type, 16#11#),
      3177 => to_slv(opcode_type, 16#17#),
      3178 => to_slv(opcode_type, 16#01#),
      3179 => to_slv(opcode_type, 16#0B#),
      3180 => to_slv(opcode_type, 16#09#),
      3181 => to_slv(opcode_type, 16#08#),
      3182 => to_slv(opcode_type, 16#03#),
      3183 => to_slv(opcode_type, 16#0C#),
      3184 => to_slv(opcode_type, 16#08#),
      3185 => to_slv(opcode_type, 16#0A#),
      3186 => to_slv(opcode_type, 16#10#),
      3187 => to_slv(opcode_type, 16#06#),
      3188 => to_slv(opcode_type, 16#07#),
      3189 => to_slv(opcode_type, 16#0F#),
      3190 => to_slv(opcode_type, 16#0A#),
      3191 => to_slv(opcode_type, 16#08#),
      3192 => to_slv(opcode_type, 16#11#),
      3193 => to_slv(opcode_type, 16#0B#),
      3194 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#09#),
      3201 => to_slv(opcode_type, 16#08#),
      3202 => to_slv(opcode_type, 16#09#),
      3203 => to_slv(opcode_type, 16#08#),
      3204 => to_slv(opcode_type, 16#0C#),
      3205 => to_slv(opcode_type, 16#0C#),
      3206 => to_slv(opcode_type, 16#09#),
      3207 => to_slv(opcode_type, 16#0B#),
      3208 => to_slv(opcode_type, 16#0D#),
      3209 => to_slv(opcode_type, 16#05#),
      3210 => to_slv(opcode_type, 16#06#),
      3211 => to_slv(opcode_type, 16#10#),
      3212 => to_slv(opcode_type, 16#0E#),
      3213 => to_slv(opcode_type, 16#06#),
      3214 => to_slv(opcode_type, 16#09#),
      3215 => to_slv(opcode_type, 16#06#),
      3216 => to_slv(opcode_type, 16#0E#),
      3217 => to_slv(opcode_type, 16#0E#),
      3218 => to_slv(opcode_type, 16#09#),
      3219 => to_slv(opcode_type, 16#10#),
      3220 => to_slv(opcode_type, 16#0C#),
      3221 => to_slv(opcode_type, 16#09#),
      3222 => to_slv(opcode_type, 16#03#),
      3223 => to_slv(opcode_type, 16#0E#),
      3224 => to_slv(opcode_type, 16#01#),
      3225 => to_slv(opcode_type, 16#0E#),
      3226 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#08#),
      3233 => to_slv(opcode_type, 16#08#),
      3234 => to_slv(opcode_type, 16#04#),
      3235 => to_slv(opcode_type, 16#03#),
      3236 => to_slv(opcode_type, 16#0D#),
      3237 => to_slv(opcode_type, 16#07#),
      3238 => to_slv(opcode_type, 16#08#),
      3239 => to_slv(opcode_type, 16#0C#),
      3240 => to_slv(opcode_type, 16#3B#),
      3241 => to_slv(opcode_type, 16#07#),
      3242 => to_slv(opcode_type, 16#0C#),
      3243 => to_slv(opcode_type, 16#0D#),
      3244 => to_slv(opcode_type, 16#09#),
      3245 => to_slv(opcode_type, 16#06#),
      3246 => to_slv(opcode_type, 16#03#),
      3247 => to_slv(opcode_type, 16#0C#),
      3248 => to_slv(opcode_type, 16#09#),
      3249 => to_slv(opcode_type, 16#5E#),
      3250 => to_slv(opcode_type, 16#0B#),
      3251 => to_slv(opcode_type, 16#07#),
      3252 => to_slv(opcode_type, 16#08#),
      3253 => to_slv(opcode_type, 16#87#),
      3254 => to_slv(opcode_type, 16#10#),
      3255 => to_slv(opcode_type, 16#08#),
      3256 => to_slv(opcode_type, 16#0B#),
      3257 => to_slv(opcode_type, 16#0B#),
      3258 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#08#),
      3265 => to_slv(opcode_type, 16#06#),
      3266 => to_slv(opcode_type, 16#08#),
      3267 => to_slv(opcode_type, 16#05#),
      3268 => to_slv(opcode_type, 16#0A#),
      3269 => to_slv(opcode_type, 16#04#),
      3270 => to_slv(opcode_type, 16#0B#),
      3271 => to_slv(opcode_type, 16#09#),
      3272 => to_slv(opcode_type, 16#01#),
      3273 => to_slv(opcode_type, 16#0E#),
      3274 => to_slv(opcode_type, 16#06#),
      3275 => to_slv(opcode_type, 16#10#),
      3276 => to_slv(opcode_type, 16#0D#),
      3277 => to_slv(opcode_type, 16#07#),
      3278 => to_slv(opcode_type, 16#06#),
      3279 => to_slv(opcode_type, 16#04#),
      3280 => to_slv(opcode_type, 16#0D#),
      3281 => to_slv(opcode_type, 16#01#),
      3282 => to_slv(opcode_type, 16#11#),
      3283 => to_slv(opcode_type, 16#07#),
      3284 => to_slv(opcode_type, 16#09#),
      3285 => to_slv(opcode_type, 16#0B#),
      3286 => to_slv(opcode_type, 16#0A#),
      3287 => to_slv(opcode_type, 16#08#),
      3288 => to_slv(opcode_type, 16#11#),
      3289 => to_slv(opcode_type, 16#0D#),
      3290 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#08#),
      3297 => to_slv(opcode_type, 16#09#),
      3298 => to_slv(opcode_type, 16#03#),
      3299 => to_slv(opcode_type, 16#09#),
      3300 => to_slv(opcode_type, 16#10#),
      3301 => to_slv(opcode_type, 16#0C#),
      3302 => to_slv(opcode_type, 16#08#),
      3303 => to_slv(opcode_type, 16#07#),
      3304 => to_slv(opcode_type, 16#10#),
      3305 => to_slv(opcode_type, 16#0F#),
      3306 => to_slv(opcode_type, 16#08#),
      3307 => to_slv(opcode_type, 16#0A#),
      3308 => to_slv(opcode_type, 16#0E#),
      3309 => to_slv(opcode_type, 16#06#),
      3310 => to_slv(opcode_type, 16#08#),
      3311 => to_slv(opcode_type, 16#06#),
      3312 => to_slv(opcode_type, 16#0C#),
      3313 => to_slv(opcode_type, 16#3C#),
      3314 => to_slv(opcode_type, 16#06#),
      3315 => to_slv(opcode_type, 16#11#),
      3316 => to_slv(opcode_type, 16#30#),
      3317 => to_slv(opcode_type, 16#08#),
      3318 => to_slv(opcode_type, 16#02#),
      3319 => to_slv(opcode_type, 16#11#),
      3320 => to_slv(opcode_type, 16#01#),
      3321 => to_slv(opcode_type, 16#C8#),
      3322 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#08#),
      3329 => to_slv(opcode_type, 16#06#),
      3330 => to_slv(opcode_type, 16#05#),
      3331 => to_slv(opcode_type, 16#05#),
      3332 => to_slv(opcode_type, 16#11#),
      3333 => to_slv(opcode_type, 16#09#),
      3334 => to_slv(opcode_type, 16#02#),
      3335 => to_slv(opcode_type, 16#0D#),
      3336 => to_slv(opcode_type, 16#08#),
      3337 => to_slv(opcode_type, 16#0D#),
      3338 => to_slv(opcode_type, 16#0D#),
      3339 => to_slv(opcode_type, 16#06#),
      3340 => to_slv(opcode_type, 16#08#),
      3341 => to_slv(opcode_type, 16#08#),
      3342 => to_slv(opcode_type, 16#0A#),
      3343 => to_slv(opcode_type, 16#0A#),
      3344 => to_slv(opcode_type, 16#07#),
      3345 => to_slv(opcode_type, 16#10#),
      3346 => to_slv(opcode_type, 16#10#),
      3347 => to_slv(opcode_type, 16#08#),
      3348 => to_slv(opcode_type, 16#09#),
      3349 => to_slv(opcode_type, 16#0F#),
      3350 => to_slv(opcode_type, 16#0B#),
      3351 => to_slv(opcode_type, 16#06#),
      3352 => to_slv(opcode_type, 16#4F#),
      3353 => to_slv(opcode_type, 16#0C#),
      3354 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#06#),
      3361 => to_slv(opcode_type, 16#06#),
      3362 => to_slv(opcode_type, 16#08#),
      3363 => to_slv(opcode_type, 16#09#),
      3364 => to_slv(opcode_type, 16#0B#),
      3365 => to_slv(opcode_type, 16#0D#),
      3366 => to_slv(opcode_type, 16#02#),
      3367 => to_slv(opcode_type, 16#0D#),
      3368 => to_slv(opcode_type, 16#07#),
      3369 => to_slv(opcode_type, 16#02#),
      3370 => to_slv(opcode_type, 16#0C#),
      3371 => to_slv(opcode_type, 16#01#),
      3372 => to_slv(opcode_type, 16#0E#),
      3373 => to_slv(opcode_type, 16#07#),
      3374 => to_slv(opcode_type, 16#08#),
      3375 => to_slv(opcode_type, 16#06#),
      3376 => to_slv(opcode_type, 16#0E#),
      3377 => to_slv(opcode_type, 16#0A#),
      3378 => to_slv(opcode_type, 16#04#),
      3379 => to_slv(opcode_type, 16#0F#),
      3380 => to_slv(opcode_type, 16#08#),
      3381 => to_slv(opcode_type, 16#09#),
      3382 => to_slv(opcode_type, 16#11#),
      3383 => to_slv(opcode_type, 16#0B#),
      3384 => to_slv(opcode_type, 16#04#),
      3385 => to_slv(opcode_type, 16#0F#),
      3386 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#09#),
      3393 => to_slv(opcode_type, 16#07#),
      3394 => to_slv(opcode_type, 16#04#),
      3395 => to_slv(opcode_type, 16#01#),
      3396 => to_slv(opcode_type, 16#0F#),
      3397 => to_slv(opcode_type, 16#06#),
      3398 => to_slv(opcode_type, 16#05#),
      3399 => to_slv(opcode_type, 16#11#),
      3400 => to_slv(opcode_type, 16#09#),
      3401 => to_slv(opcode_type, 16#0A#),
      3402 => to_slv(opcode_type, 16#0B#),
      3403 => to_slv(opcode_type, 16#09#),
      3404 => to_slv(opcode_type, 16#07#),
      3405 => to_slv(opcode_type, 16#08#),
      3406 => to_slv(opcode_type, 16#0E#),
      3407 => to_slv(opcode_type, 16#11#),
      3408 => to_slv(opcode_type, 16#06#),
      3409 => to_slv(opcode_type, 16#0E#),
      3410 => to_slv(opcode_type, 16#0E#),
      3411 => to_slv(opcode_type, 16#07#),
      3412 => to_slv(opcode_type, 16#09#),
      3413 => to_slv(opcode_type, 16#11#),
      3414 => to_slv(opcode_type, 16#BF#),
      3415 => to_slv(opcode_type, 16#06#),
      3416 => to_slv(opcode_type, 16#2F#),
      3417 => to_slv(opcode_type, 16#0D#),
      3418 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#07#),
      3425 => to_slv(opcode_type, 16#07#),
      3426 => to_slv(opcode_type, 16#03#),
      3427 => to_slv(opcode_type, 16#09#),
      3428 => to_slv(opcode_type, 16#0E#),
      3429 => to_slv(opcode_type, 16#0F#),
      3430 => to_slv(opcode_type, 16#07#),
      3431 => to_slv(opcode_type, 16#05#),
      3432 => to_slv(opcode_type, 16#54#),
      3433 => to_slv(opcode_type, 16#04#),
      3434 => to_slv(opcode_type, 16#0A#),
      3435 => to_slv(opcode_type, 16#06#),
      3436 => to_slv(opcode_type, 16#09#),
      3437 => to_slv(opcode_type, 16#06#),
      3438 => to_slv(opcode_type, 16#0D#),
      3439 => to_slv(opcode_type, 16#0B#),
      3440 => to_slv(opcode_type, 16#07#),
      3441 => to_slv(opcode_type, 16#E7#),
      3442 => to_slv(opcode_type, 16#10#),
      3443 => to_slv(opcode_type, 16#06#),
      3444 => to_slv(opcode_type, 16#09#),
      3445 => to_slv(opcode_type, 16#0C#),
      3446 => to_slv(opcode_type, 16#0C#),
      3447 => to_slv(opcode_type, 16#08#),
      3448 => to_slv(opcode_type, 16#0B#),
      3449 => to_slv(opcode_type, 16#0E#),
      3450 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#07#),
      3457 => to_slv(opcode_type, 16#08#),
      3458 => to_slv(opcode_type, 16#09#),
      3459 => to_slv(opcode_type, 16#04#),
      3460 => to_slv(opcode_type, 16#0E#),
      3461 => to_slv(opcode_type, 16#05#),
      3462 => to_slv(opcode_type, 16#0E#),
      3463 => to_slv(opcode_type, 16#07#),
      3464 => to_slv(opcode_type, 16#06#),
      3465 => to_slv(opcode_type, 16#0E#),
      3466 => to_slv(opcode_type, 16#0C#),
      3467 => to_slv(opcode_type, 16#08#),
      3468 => to_slv(opcode_type, 16#7C#),
      3469 => to_slv(opcode_type, 16#0C#),
      3470 => to_slv(opcode_type, 16#08#),
      3471 => to_slv(opcode_type, 16#01#),
      3472 => to_slv(opcode_type, 16#07#),
      3473 => to_slv(opcode_type, 16#0B#),
      3474 => to_slv(opcode_type, 16#10#),
      3475 => to_slv(opcode_type, 16#08#),
      3476 => to_slv(opcode_type, 16#07#),
      3477 => to_slv(opcode_type, 16#0B#),
      3478 => to_slv(opcode_type, 16#0B#),
      3479 => to_slv(opcode_type, 16#09#),
      3480 => to_slv(opcode_type, 16#0C#),
      3481 => to_slv(opcode_type, 16#0F#),
      3482 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#08#),
      3489 => to_slv(opcode_type, 16#07#),
      3490 => to_slv(opcode_type, 16#04#),
      3491 => to_slv(opcode_type, 16#05#),
      3492 => to_slv(opcode_type, 16#10#),
      3493 => to_slv(opcode_type, 16#06#),
      3494 => to_slv(opcode_type, 16#04#),
      3495 => to_slv(opcode_type, 16#11#),
      3496 => to_slv(opcode_type, 16#09#),
      3497 => to_slv(opcode_type, 16#6F#),
      3498 => to_slv(opcode_type, 16#0A#),
      3499 => to_slv(opcode_type, 16#06#),
      3500 => to_slv(opcode_type, 16#07#),
      3501 => to_slv(opcode_type, 16#09#),
      3502 => to_slv(opcode_type, 16#0D#),
      3503 => to_slv(opcode_type, 16#0C#),
      3504 => to_slv(opcode_type, 16#07#),
      3505 => to_slv(opcode_type, 16#11#),
      3506 => to_slv(opcode_type, 16#11#),
      3507 => to_slv(opcode_type, 16#09#),
      3508 => to_slv(opcode_type, 16#08#),
      3509 => to_slv(opcode_type, 16#76#),
      3510 => to_slv(opcode_type, 16#11#),
      3511 => to_slv(opcode_type, 16#06#),
      3512 => to_slv(opcode_type, 16#90#),
      3513 => to_slv(opcode_type, 16#0E#),
      3514 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#09#),
      3521 => to_slv(opcode_type, 16#09#),
      3522 => to_slv(opcode_type, 16#05#),
      3523 => to_slv(opcode_type, 16#09#),
      3524 => to_slv(opcode_type, 16#0B#),
      3525 => to_slv(opcode_type, 16#0D#),
      3526 => to_slv(opcode_type, 16#06#),
      3527 => to_slv(opcode_type, 16#08#),
      3528 => to_slv(opcode_type, 16#0B#),
      3529 => to_slv(opcode_type, 16#0C#),
      3530 => to_slv(opcode_type, 16#07#),
      3531 => to_slv(opcode_type, 16#11#),
      3532 => to_slv(opcode_type, 16#D7#),
      3533 => to_slv(opcode_type, 16#06#),
      3534 => to_slv(opcode_type, 16#08#),
      3535 => to_slv(opcode_type, 16#01#),
      3536 => to_slv(opcode_type, 16#0E#),
      3537 => to_slv(opcode_type, 16#09#),
      3538 => to_slv(opcode_type, 16#28#),
      3539 => to_slv(opcode_type, 16#0E#),
      3540 => to_slv(opcode_type, 16#06#),
      3541 => to_slv(opcode_type, 16#09#),
      3542 => to_slv(opcode_type, 16#11#),
      3543 => to_slv(opcode_type, 16#10#),
      3544 => to_slv(opcode_type, 16#04#),
      3545 => to_slv(opcode_type, 16#0A#),
      3546 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#08#),
      3553 => to_slv(opcode_type, 16#06#),
      3554 => to_slv(opcode_type, 16#04#),
      3555 => to_slv(opcode_type, 16#04#),
      3556 => to_slv(opcode_type, 16#10#),
      3557 => to_slv(opcode_type, 16#09#),
      3558 => to_slv(opcode_type, 16#05#),
      3559 => to_slv(opcode_type, 16#0B#),
      3560 => to_slv(opcode_type, 16#07#),
      3561 => to_slv(opcode_type, 16#0F#),
      3562 => to_slv(opcode_type, 16#0B#),
      3563 => to_slv(opcode_type, 16#09#),
      3564 => to_slv(opcode_type, 16#06#),
      3565 => to_slv(opcode_type, 16#06#),
      3566 => to_slv(opcode_type, 16#0C#),
      3567 => to_slv(opcode_type, 16#0D#),
      3568 => to_slv(opcode_type, 16#08#),
      3569 => to_slv(opcode_type, 16#C4#),
      3570 => to_slv(opcode_type, 16#10#),
      3571 => to_slv(opcode_type, 16#08#),
      3572 => to_slv(opcode_type, 16#09#),
      3573 => to_slv(opcode_type, 16#0A#),
      3574 => to_slv(opcode_type, 16#0E#),
      3575 => to_slv(opcode_type, 16#06#),
      3576 => to_slv(opcode_type, 16#0C#),
      3577 => to_slv(opcode_type, 16#0D#),
      3578 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#07#),
      3585 => to_slv(opcode_type, 16#06#),
      3586 => to_slv(opcode_type, 16#08#),
      3587 => to_slv(opcode_type, 16#05#),
      3588 => to_slv(opcode_type, 16#1F#),
      3589 => to_slv(opcode_type, 16#02#),
      3590 => to_slv(opcode_type, 16#0E#),
      3591 => to_slv(opcode_type, 16#09#),
      3592 => to_slv(opcode_type, 16#05#),
      3593 => to_slv(opcode_type, 16#11#),
      3594 => to_slv(opcode_type, 16#07#),
      3595 => to_slv(opcode_type, 16#10#),
      3596 => to_slv(opcode_type, 16#0D#),
      3597 => to_slv(opcode_type, 16#08#),
      3598 => to_slv(opcode_type, 16#07#),
      3599 => to_slv(opcode_type, 16#06#),
      3600 => to_slv(opcode_type, 16#0B#),
      3601 => to_slv(opcode_type, 16#10#),
      3602 => to_slv(opcode_type, 16#04#),
      3603 => to_slv(opcode_type, 16#0D#),
      3604 => to_slv(opcode_type, 16#06#),
      3605 => to_slv(opcode_type, 16#03#),
      3606 => to_slv(opcode_type, 16#11#),
      3607 => to_slv(opcode_type, 16#08#),
      3608 => to_slv(opcode_type, 16#0E#),
      3609 => to_slv(opcode_type, 16#0B#),
      3610 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#07#),
      3617 => to_slv(opcode_type, 16#09#),
      3618 => to_slv(opcode_type, 16#04#),
      3619 => to_slv(opcode_type, 16#02#),
      3620 => to_slv(opcode_type, 16#9C#),
      3621 => to_slv(opcode_type, 16#07#),
      3622 => to_slv(opcode_type, 16#08#),
      3623 => to_slv(opcode_type, 16#0C#),
      3624 => to_slv(opcode_type, 16#0D#),
      3625 => to_slv(opcode_type, 16#01#),
      3626 => to_slv(opcode_type, 16#0F#),
      3627 => to_slv(opcode_type, 16#07#),
      3628 => to_slv(opcode_type, 16#08#),
      3629 => to_slv(opcode_type, 16#09#),
      3630 => to_slv(opcode_type, 16#0B#),
      3631 => to_slv(opcode_type, 16#11#),
      3632 => to_slv(opcode_type, 16#06#),
      3633 => to_slv(opcode_type, 16#10#),
      3634 => to_slv(opcode_type, 16#0E#),
      3635 => to_slv(opcode_type, 16#07#),
      3636 => to_slv(opcode_type, 16#07#),
      3637 => to_slv(opcode_type, 16#11#),
      3638 => to_slv(opcode_type, 16#11#),
      3639 => to_slv(opcode_type, 16#07#),
      3640 => to_slv(opcode_type, 16#0C#),
      3641 => to_slv(opcode_type, 16#11#),
      3642 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#08#),
      3649 => to_slv(opcode_type, 16#06#),
      3650 => to_slv(opcode_type, 16#06#),
      3651 => to_slv(opcode_type, 16#04#),
      3652 => to_slv(opcode_type, 16#0F#),
      3653 => to_slv(opcode_type, 16#03#),
      3654 => to_slv(opcode_type, 16#0C#),
      3655 => to_slv(opcode_type, 16#06#),
      3656 => to_slv(opcode_type, 16#06#),
      3657 => to_slv(opcode_type, 16#0C#),
      3658 => to_slv(opcode_type, 16#0B#),
      3659 => to_slv(opcode_type, 16#09#),
      3660 => to_slv(opcode_type, 16#0F#),
      3661 => to_slv(opcode_type, 16#0B#),
      3662 => to_slv(opcode_type, 16#07#),
      3663 => to_slv(opcode_type, 16#01#),
      3664 => to_slv(opcode_type, 16#06#),
      3665 => to_slv(opcode_type, 16#0C#),
      3666 => to_slv(opcode_type, 16#0E#),
      3667 => to_slv(opcode_type, 16#08#),
      3668 => to_slv(opcode_type, 16#08#),
      3669 => to_slv(opcode_type, 16#F7#),
      3670 => to_slv(opcode_type, 16#10#),
      3671 => to_slv(opcode_type, 16#09#),
      3672 => to_slv(opcode_type, 16#0E#),
      3673 => to_slv(opcode_type, 16#0D#),
      3674 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#06#),
      3681 => to_slv(opcode_type, 16#06#),
      3682 => to_slv(opcode_type, 16#07#),
      3683 => to_slv(opcode_type, 16#06#),
      3684 => to_slv(opcode_type, 16#0C#),
      3685 => to_slv(opcode_type, 16#0D#),
      3686 => to_slv(opcode_type, 16#01#),
      3687 => to_slv(opcode_type, 16#0C#),
      3688 => to_slv(opcode_type, 16#08#),
      3689 => to_slv(opcode_type, 16#03#),
      3690 => to_slv(opcode_type, 16#0D#),
      3691 => to_slv(opcode_type, 16#02#),
      3692 => to_slv(opcode_type, 16#0E#),
      3693 => to_slv(opcode_type, 16#08#),
      3694 => to_slv(opcode_type, 16#07#),
      3695 => to_slv(opcode_type, 16#05#),
      3696 => to_slv(opcode_type, 16#0E#),
      3697 => to_slv(opcode_type, 16#08#),
      3698 => to_slv(opcode_type, 16#10#),
      3699 => to_slv(opcode_type, 16#0E#),
      3700 => to_slv(opcode_type, 16#09#),
      3701 => to_slv(opcode_type, 16#05#),
      3702 => to_slv(opcode_type, 16#10#),
      3703 => to_slv(opcode_type, 16#06#),
      3704 => to_slv(opcode_type, 16#0B#),
      3705 => to_slv(opcode_type, 16#11#),
      3706 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#07#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#08#),
      3715 => to_slv(opcode_type, 16#05#),
      3716 => to_slv(opcode_type, 16#0D#),
      3717 => to_slv(opcode_type, 16#06#),
      3718 => to_slv(opcode_type, 16#0F#),
      3719 => to_slv(opcode_type, 16#10#),
      3720 => to_slv(opcode_type, 16#04#),
      3721 => to_slv(opcode_type, 16#03#),
      3722 => to_slv(opcode_type, 16#0A#),
      3723 => to_slv(opcode_type, 16#07#),
      3724 => to_slv(opcode_type, 16#06#),
      3725 => to_slv(opcode_type, 16#06#),
      3726 => to_slv(opcode_type, 16#10#),
      3727 => to_slv(opcode_type, 16#0E#),
      3728 => to_slv(opcode_type, 16#09#),
      3729 => to_slv(opcode_type, 16#0B#),
      3730 => to_slv(opcode_type, 16#0F#),
      3731 => to_slv(opcode_type, 16#08#),
      3732 => to_slv(opcode_type, 16#07#),
      3733 => to_slv(opcode_type, 16#11#),
      3734 => to_slv(opcode_type, 16#0D#),
      3735 => to_slv(opcode_type, 16#09#),
      3736 => to_slv(opcode_type, 16#10#),
      3737 => to_slv(opcode_type, 16#0F#),
      3738 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#09#),
      3745 => to_slv(opcode_type, 16#09#),
      3746 => to_slv(opcode_type, 16#03#),
      3747 => to_slv(opcode_type, 16#07#),
      3748 => to_slv(opcode_type, 16#0E#),
      3749 => to_slv(opcode_type, 16#0C#),
      3750 => to_slv(opcode_type, 16#08#),
      3751 => to_slv(opcode_type, 16#06#),
      3752 => to_slv(opcode_type, 16#0C#),
      3753 => to_slv(opcode_type, 16#0D#),
      3754 => to_slv(opcode_type, 16#02#),
      3755 => to_slv(opcode_type, 16#10#),
      3756 => to_slv(opcode_type, 16#09#),
      3757 => to_slv(opcode_type, 16#09#),
      3758 => to_slv(opcode_type, 16#04#),
      3759 => to_slv(opcode_type, 16#11#),
      3760 => to_slv(opcode_type, 16#09#),
      3761 => to_slv(opcode_type, 16#0A#),
      3762 => to_slv(opcode_type, 16#11#),
      3763 => to_slv(opcode_type, 16#06#),
      3764 => to_slv(opcode_type, 16#06#),
      3765 => to_slv(opcode_type, 16#68#),
      3766 => to_slv(opcode_type, 16#0A#),
      3767 => to_slv(opcode_type, 16#09#),
      3768 => to_slv(opcode_type, 16#10#),
      3769 => to_slv(opcode_type, 16#0E#),
      3770 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#07#),
      3777 => to_slv(opcode_type, 16#07#),
      3778 => to_slv(opcode_type, 16#06#),
      3779 => to_slv(opcode_type, 16#07#),
      3780 => to_slv(opcode_type, 16#10#),
      3781 => to_slv(opcode_type, 16#0F#),
      3782 => to_slv(opcode_type, 16#09#),
      3783 => to_slv(opcode_type, 16#11#),
      3784 => to_slv(opcode_type, 16#0E#),
      3785 => to_slv(opcode_type, 16#06#),
      3786 => to_slv(opcode_type, 16#05#),
      3787 => to_slv(opcode_type, 16#10#),
      3788 => to_slv(opcode_type, 16#09#),
      3789 => to_slv(opcode_type, 16#0C#),
      3790 => to_slv(opcode_type, 16#0D#),
      3791 => to_slv(opcode_type, 16#08#),
      3792 => to_slv(opcode_type, 16#05#),
      3793 => to_slv(opcode_type, 16#02#),
      3794 => to_slv(opcode_type, 16#11#),
      3795 => to_slv(opcode_type, 16#09#),
      3796 => to_slv(opcode_type, 16#07#),
      3797 => to_slv(opcode_type, 16#0F#),
      3798 => to_slv(opcode_type, 16#0F#),
      3799 => to_slv(opcode_type, 16#08#),
      3800 => to_slv(opcode_type, 16#0A#),
      3801 => to_slv(opcode_type, 16#0E#),
      3802 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#08#),
      3809 => to_slv(opcode_type, 16#07#),
      3810 => to_slv(opcode_type, 16#01#),
      3811 => to_slv(opcode_type, 16#06#),
      3812 => to_slv(opcode_type, 16#66#),
      3813 => to_slv(opcode_type, 16#0F#),
      3814 => to_slv(opcode_type, 16#09#),
      3815 => to_slv(opcode_type, 16#06#),
      3816 => to_slv(opcode_type, 16#0D#),
      3817 => to_slv(opcode_type, 16#0C#),
      3818 => to_slv(opcode_type, 16#06#),
      3819 => to_slv(opcode_type, 16#10#),
      3820 => to_slv(opcode_type, 16#0A#),
      3821 => to_slv(opcode_type, 16#07#),
      3822 => to_slv(opcode_type, 16#07#),
      3823 => to_slv(opcode_type, 16#04#),
      3824 => to_slv(opcode_type, 16#0B#),
      3825 => to_slv(opcode_type, 16#05#),
      3826 => to_slv(opcode_type, 16#0A#),
      3827 => to_slv(opcode_type, 16#06#),
      3828 => to_slv(opcode_type, 16#09#),
      3829 => to_slv(opcode_type, 16#0D#),
      3830 => to_slv(opcode_type, 16#0F#),
      3831 => to_slv(opcode_type, 16#08#),
      3832 => to_slv(opcode_type, 16#0D#),
      3833 => to_slv(opcode_type, 16#10#),
      3834 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#06#),
      3841 => to_slv(opcode_type, 16#09#),
      3842 => to_slv(opcode_type, 16#01#),
      3843 => to_slv(opcode_type, 16#01#),
      3844 => to_slv(opcode_type, 16#0E#),
      3845 => to_slv(opcode_type, 16#08#),
      3846 => to_slv(opcode_type, 16#01#),
      3847 => to_slv(opcode_type, 16#27#),
      3848 => to_slv(opcode_type, 16#07#),
      3849 => to_slv(opcode_type, 16#0C#),
      3850 => to_slv(opcode_type, 16#10#),
      3851 => to_slv(opcode_type, 16#06#),
      3852 => to_slv(opcode_type, 16#07#),
      3853 => to_slv(opcode_type, 16#07#),
      3854 => to_slv(opcode_type, 16#0F#),
      3855 => to_slv(opcode_type, 16#10#),
      3856 => to_slv(opcode_type, 16#08#),
      3857 => to_slv(opcode_type, 16#0A#),
      3858 => to_slv(opcode_type, 16#0A#),
      3859 => to_slv(opcode_type, 16#06#),
      3860 => to_slv(opcode_type, 16#07#),
      3861 => to_slv(opcode_type, 16#0D#),
      3862 => to_slv(opcode_type, 16#7E#),
      3863 => to_slv(opcode_type, 16#06#),
      3864 => to_slv(opcode_type, 16#0D#),
      3865 => to_slv(opcode_type, 16#11#),
      3866 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#08#),
      3873 => to_slv(opcode_type, 16#09#),
      3874 => to_slv(opcode_type, 16#06#),
      3875 => to_slv(opcode_type, 16#07#),
      3876 => to_slv(opcode_type, 16#0C#),
      3877 => to_slv(opcode_type, 16#0F#),
      3878 => to_slv(opcode_type, 16#07#),
      3879 => to_slv(opcode_type, 16#0D#),
      3880 => to_slv(opcode_type, 16#71#),
      3881 => to_slv(opcode_type, 16#08#),
      3882 => to_slv(opcode_type, 16#08#),
      3883 => to_slv(opcode_type, 16#10#),
      3884 => to_slv(opcode_type, 16#10#),
      3885 => to_slv(opcode_type, 16#06#),
      3886 => to_slv(opcode_type, 16#0A#),
      3887 => to_slv(opcode_type, 16#0C#),
      3888 => to_slv(opcode_type, 16#09#),
      3889 => to_slv(opcode_type, 16#09#),
      3890 => to_slv(opcode_type, 16#02#),
      3891 => to_slv(opcode_type, 16#0F#),
      3892 => to_slv(opcode_type, 16#01#),
      3893 => to_slv(opcode_type, 16#11#),
      3894 => to_slv(opcode_type, 16#02#),
      3895 => to_slv(opcode_type, 16#06#),
      3896 => to_slv(opcode_type, 16#0F#),
      3897 => to_slv(opcode_type, 16#0E#),
      3898 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#06#),
      3905 => to_slv(opcode_type, 16#07#),
      3906 => to_slv(opcode_type, 16#04#),
      3907 => to_slv(opcode_type, 16#09#),
      3908 => to_slv(opcode_type, 16#CB#),
      3909 => to_slv(opcode_type, 16#10#),
      3910 => to_slv(opcode_type, 16#07#),
      3911 => to_slv(opcode_type, 16#09#),
      3912 => to_slv(opcode_type, 16#0B#),
      3913 => to_slv(opcode_type, 16#0B#),
      3914 => to_slv(opcode_type, 16#04#),
      3915 => to_slv(opcode_type, 16#0D#),
      3916 => to_slv(opcode_type, 16#07#),
      3917 => to_slv(opcode_type, 16#07#),
      3918 => to_slv(opcode_type, 16#01#),
      3919 => to_slv(opcode_type, 16#0E#),
      3920 => to_slv(opcode_type, 16#06#),
      3921 => to_slv(opcode_type, 16#0F#),
      3922 => to_slv(opcode_type, 16#0E#),
      3923 => to_slv(opcode_type, 16#06#),
      3924 => to_slv(opcode_type, 16#09#),
      3925 => to_slv(opcode_type, 16#0D#),
      3926 => to_slv(opcode_type, 16#11#),
      3927 => to_slv(opcode_type, 16#09#),
      3928 => to_slv(opcode_type, 16#0D#),
      3929 => to_slv(opcode_type, 16#11#),
      3930 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#06#),
      3937 => to_slv(opcode_type, 16#09#),
      3938 => to_slv(opcode_type, 16#04#),
      3939 => to_slv(opcode_type, 16#05#),
      3940 => to_slv(opcode_type, 16#0D#),
      3941 => to_slv(opcode_type, 16#07#),
      3942 => to_slv(opcode_type, 16#01#),
      3943 => to_slv(opcode_type, 16#0A#),
      3944 => to_slv(opcode_type, 16#08#),
      3945 => to_slv(opcode_type, 16#11#),
      3946 => to_slv(opcode_type, 16#11#),
      3947 => to_slv(opcode_type, 16#06#),
      3948 => to_slv(opcode_type, 16#08#),
      3949 => to_slv(opcode_type, 16#07#),
      3950 => to_slv(opcode_type, 16#0E#),
      3951 => to_slv(opcode_type, 16#0A#),
      3952 => to_slv(opcode_type, 16#09#),
      3953 => to_slv(opcode_type, 16#8C#),
      3954 => to_slv(opcode_type, 16#0A#),
      3955 => to_slv(opcode_type, 16#07#),
      3956 => to_slv(opcode_type, 16#08#),
      3957 => to_slv(opcode_type, 16#11#),
      3958 => to_slv(opcode_type, 16#10#),
      3959 => to_slv(opcode_type, 16#09#),
      3960 => to_slv(opcode_type, 16#0F#),
      3961 => to_slv(opcode_type, 16#0E#),
      3962 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#08#),
      3969 => to_slv(opcode_type, 16#07#),
      3970 => to_slv(opcode_type, 16#08#),
      3971 => to_slv(opcode_type, 16#09#),
      3972 => to_slv(opcode_type, 16#0E#),
      3973 => to_slv(opcode_type, 16#0A#),
      3974 => to_slv(opcode_type, 16#04#),
      3975 => to_slv(opcode_type, 16#77#),
      3976 => to_slv(opcode_type, 16#04#),
      3977 => to_slv(opcode_type, 16#02#),
      3978 => to_slv(opcode_type, 16#0D#),
      3979 => to_slv(opcode_type, 16#09#),
      3980 => to_slv(opcode_type, 16#06#),
      3981 => to_slv(opcode_type, 16#07#),
      3982 => to_slv(opcode_type, 16#0D#),
      3983 => to_slv(opcode_type, 16#0F#),
      3984 => to_slv(opcode_type, 16#06#),
      3985 => to_slv(opcode_type, 16#0D#),
      3986 => to_slv(opcode_type, 16#11#),
      3987 => to_slv(opcode_type, 16#06#),
      3988 => to_slv(opcode_type, 16#06#),
      3989 => to_slv(opcode_type, 16#0B#),
      3990 => to_slv(opcode_type, 16#0B#),
      3991 => to_slv(opcode_type, 16#06#),
      3992 => to_slv(opcode_type, 16#0E#),
      3993 => to_slv(opcode_type, 16#0E#),
      3994 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#07#),
      4001 => to_slv(opcode_type, 16#06#),
      4002 => to_slv(opcode_type, 16#09#),
      4003 => to_slv(opcode_type, 16#05#),
      4004 => to_slv(opcode_type, 16#0D#),
      4005 => to_slv(opcode_type, 16#01#),
      4006 => to_slv(opcode_type, 16#0D#),
      4007 => to_slv(opcode_type, 16#07#),
      4008 => to_slv(opcode_type, 16#06#),
      4009 => to_slv(opcode_type, 16#0E#),
      4010 => to_slv(opcode_type, 16#0D#),
      4011 => to_slv(opcode_type, 16#06#),
      4012 => to_slv(opcode_type, 16#10#),
      4013 => to_slv(opcode_type, 16#0B#),
      4014 => to_slv(opcode_type, 16#09#),
      4015 => to_slv(opcode_type, 16#06#),
      4016 => to_slv(opcode_type, 16#04#),
      4017 => to_slv(opcode_type, 16#0B#),
      4018 => to_slv(opcode_type, 16#06#),
      4019 => to_slv(opcode_type, 16#22#),
      4020 => to_slv(opcode_type, 16#0C#),
      4021 => to_slv(opcode_type, 16#07#),
      4022 => to_slv(opcode_type, 16#04#),
      4023 => to_slv(opcode_type, 16#0D#),
      4024 => to_slv(opcode_type, 16#01#),
      4025 => to_slv(opcode_type, 16#0C#),
      4026 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#08#),
      4033 => to_slv(opcode_type, 16#06#),
      4034 => to_slv(opcode_type, 16#05#),
      4035 => to_slv(opcode_type, 16#07#),
      4036 => to_slv(opcode_type, 16#2F#),
      4037 => to_slv(opcode_type, 16#7F#),
      4038 => to_slv(opcode_type, 16#06#),
      4039 => to_slv(opcode_type, 16#04#),
      4040 => to_slv(opcode_type, 16#0D#),
      4041 => to_slv(opcode_type, 16#07#),
      4042 => to_slv(opcode_type, 16#0A#),
      4043 => to_slv(opcode_type, 16#10#),
      4044 => to_slv(opcode_type, 16#09#),
      4045 => to_slv(opcode_type, 16#08#),
      4046 => to_slv(opcode_type, 16#09#),
      4047 => to_slv(opcode_type, 16#0B#),
      4048 => to_slv(opcode_type, 16#10#),
      4049 => to_slv(opcode_type, 16#08#),
      4050 => to_slv(opcode_type, 16#0B#),
      4051 => to_slv(opcode_type, 16#0F#),
      4052 => to_slv(opcode_type, 16#09#),
      4053 => to_slv(opcode_type, 16#07#),
      4054 => to_slv(opcode_type, 16#BE#),
      4055 => to_slv(opcode_type, 16#0E#),
      4056 => to_slv(opcode_type, 16#02#),
      4057 => to_slv(opcode_type, 16#0B#),
      4058 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#08#),
      4066 => to_slv(opcode_type, 16#08#),
      4067 => to_slv(opcode_type, 16#08#),
      4068 => to_slv(opcode_type, 16#0C#),
      4069 => to_slv(opcode_type, 16#11#),
      4070 => to_slv(opcode_type, 16#03#),
      4071 => to_slv(opcode_type, 16#E3#),
      4072 => to_slv(opcode_type, 16#03#),
      4073 => to_slv(opcode_type, 16#04#),
      4074 => to_slv(opcode_type, 16#11#),
      4075 => to_slv(opcode_type, 16#09#),
      4076 => to_slv(opcode_type, 16#08#),
      4077 => to_slv(opcode_type, 16#08#),
      4078 => to_slv(opcode_type, 16#0B#),
      4079 => to_slv(opcode_type, 16#0D#),
      4080 => to_slv(opcode_type, 16#07#),
      4081 => to_slv(opcode_type, 16#0D#),
      4082 => to_slv(opcode_type, 16#10#),
      4083 => to_slv(opcode_type, 16#08#),
      4084 => to_slv(opcode_type, 16#07#),
      4085 => to_slv(opcode_type, 16#10#),
      4086 => to_slv(opcode_type, 16#0C#),
      4087 => to_slv(opcode_type, 16#06#),
      4088 => to_slv(opcode_type, 16#0A#),
      4089 => to_slv(opcode_type, 16#0B#),
      4090 to 4095 => (others => '0')
  ),

    -- Bin `27`...
    26 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#07#),
      1 => to_slv(opcode_type, 16#09#),
      2 => to_slv(opcode_type, 16#01#),
      3 => to_slv(opcode_type, 16#01#),
      4 => to_slv(opcode_type, 16#0F#),
      5 => to_slv(opcode_type, 16#06#),
      6 => to_slv(opcode_type, 16#09#),
      7 => to_slv(opcode_type, 16#10#),
      8 => to_slv(opcode_type, 16#10#),
      9 => to_slv(opcode_type, 16#08#),
      10 => to_slv(opcode_type, 16#11#),
      11 => to_slv(opcode_type, 16#11#),
      12 => to_slv(opcode_type, 16#06#),
      13 => to_slv(opcode_type, 16#08#),
      14 => to_slv(opcode_type, 16#07#),
      15 => to_slv(opcode_type, 16#11#),
      16 => to_slv(opcode_type, 16#11#),
      17 => to_slv(opcode_type, 16#09#),
      18 => to_slv(opcode_type, 16#0F#),
      19 => to_slv(opcode_type, 16#0D#),
      20 => to_slv(opcode_type, 16#08#),
      21 => to_slv(opcode_type, 16#07#),
      22 => to_slv(opcode_type, 16#28#),
      23 => to_slv(opcode_type, 16#0F#),
      24 => to_slv(opcode_type, 16#07#),
      25 => to_slv(opcode_type, 16#0A#),
      26 => to_slv(opcode_type, 16#0E#),
      27 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#08#),
      33 => to_slv(opcode_type, 16#09#),
      34 => to_slv(opcode_type, 16#05#),
      35 => to_slv(opcode_type, 16#07#),
      36 => to_slv(opcode_type, 16#10#),
      37 => to_slv(opcode_type, 16#0D#),
      38 => to_slv(opcode_type, 16#08#),
      39 => to_slv(opcode_type, 16#08#),
      40 => to_slv(opcode_type, 16#E0#),
      41 => to_slv(opcode_type, 16#11#),
      42 => to_slv(opcode_type, 16#07#),
      43 => to_slv(opcode_type, 16#0D#),
      44 => to_slv(opcode_type, 16#0E#),
      45 => to_slv(opcode_type, 16#07#),
      46 => to_slv(opcode_type, 16#07#),
      47 => to_slv(opcode_type, 16#06#),
      48 => to_slv(opcode_type, 16#0D#),
      49 => to_slv(opcode_type, 16#0E#),
      50 => to_slv(opcode_type, 16#05#),
      51 => to_slv(opcode_type, 16#10#),
      52 => to_slv(opcode_type, 16#06#),
      53 => to_slv(opcode_type, 16#08#),
      54 => to_slv(opcode_type, 16#0A#),
      55 => to_slv(opcode_type, 16#10#),
      56 => to_slv(opcode_type, 16#08#),
      57 => to_slv(opcode_type, 16#0F#),
      58 => to_slv(opcode_type, 16#0F#),
      59 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#06#),
      65 => to_slv(opcode_type, 16#06#),
      66 => to_slv(opcode_type, 16#02#),
      67 => to_slv(opcode_type, 16#09#),
      68 => to_slv(opcode_type, 16#BB#),
      69 => to_slv(opcode_type, 16#AE#),
      70 => to_slv(opcode_type, 16#09#),
      71 => to_slv(opcode_type, 16#02#),
      72 => to_slv(opcode_type, 16#0D#),
      73 => to_slv(opcode_type, 16#07#),
      74 => to_slv(opcode_type, 16#11#),
      75 => to_slv(opcode_type, 16#10#),
      76 => to_slv(opcode_type, 16#07#),
      77 => to_slv(opcode_type, 16#07#),
      78 => to_slv(opcode_type, 16#06#),
      79 => to_slv(opcode_type, 16#10#),
      80 => to_slv(opcode_type, 16#0F#),
      81 => to_slv(opcode_type, 16#07#),
      82 => to_slv(opcode_type, 16#0B#),
      83 => to_slv(opcode_type, 16#11#),
      84 => to_slv(opcode_type, 16#09#),
      85 => to_slv(opcode_type, 16#07#),
      86 => to_slv(opcode_type, 16#0D#),
      87 => to_slv(opcode_type, 16#89#),
      88 => to_slv(opcode_type, 16#07#),
      89 => to_slv(opcode_type, 16#10#),
      90 => to_slv(opcode_type, 16#11#),
      91 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#09#),
      97 => to_slv(opcode_type, 16#08#),
      98 => to_slv(opcode_type, 16#02#),
      99 => to_slv(opcode_type, 16#04#),
      100 => to_slv(opcode_type, 16#BA#),
      101 => to_slv(opcode_type, 16#07#),
      102 => to_slv(opcode_type, 16#06#),
      103 => to_slv(opcode_type, 16#10#),
      104 => to_slv(opcode_type, 16#10#),
      105 => to_slv(opcode_type, 16#08#),
      106 => to_slv(opcode_type, 16#0E#),
      107 => to_slv(opcode_type, 16#0F#),
      108 => to_slv(opcode_type, 16#06#),
      109 => to_slv(opcode_type, 16#06#),
      110 => to_slv(opcode_type, 16#06#),
      111 => to_slv(opcode_type, 16#0A#),
      112 => to_slv(opcode_type, 16#0C#),
      113 => to_slv(opcode_type, 16#07#),
      114 => to_slv(opcode_type, 16#0D#),
      115 => to_slv(opcode_type, 16#D2#),
      116 => to_slv(opcode_type, 16#07#),
      117 => to_slv(opcode_type, 16#09#),
      118 => to_slv(opcode_type, 16#0B#),
      119 => to_slv(opcode_type, 16#11#),
      120 => to_slv(opcode_type, 16#09#),
      121 => to_slv(opcode_type, 16#E6#),
      122 => to_slv(opcode_type, 16#0F#),
      123 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#09#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#04#),
      131 => to_slv(opcode_type, 16#08#),
      132 => to_slv(opcode_type, 16#0C#),
      133 => to_slv(opcode_type, 16#0B#),
      134 => to_slv(opcode_type, 16#09#),
      135 => to_slv(opcode_type, 16#01#),
      136 => to_slv(opcode_type, 16#10#),
      137 => to_slv(opcode_type, 16#07#),
      138 => to_slv(opcode_type, 16#0D#),
      139 => to_slv(opcode_type, 16#0B#),
      140 => to_slv(opcode_type, 16#06#),
      141 => to_slv(opcode_type, 16#07#),
      142 => to_slv(opcode_type, 16#09#),
      143 => to_slv(opcode_type, 16#19#),
      144 => to_slv(opcode_type, 16#11#),
      145 => to_slv(opcode_type, 16#09#),
      146 => to_slv(opcode_type, 16#0D#),
      147 => to_slv(opcode_type, 16#0C#),
      148 => to_slv(opcode_type, 16#08#),
      149 => to_slv(opcode_type, 16#06#),
      150 => to_slv(opcode_type, 16#0F#),
      151 => to_slv(opcode_type, 16#0C#),
      152 => to_slv(opcode_type, 16#06#),
      153 => to_slv(opcode_type, 16#11#),
      154 => to_slv(opcode_type, 16#11#),
      155 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#07#),
      161 => to_slv(opcode_type, 16#09#),
      162 => to_slv(opcode_type, 16#01#),
      163 => to_slv(opcode_type, 16#07#),
      164 => to_slv(opcode_type, 16#0C#),
      165 => to_slv(opcode_type, 16#0D#),
      166 => to_slv(opcode_type, 16#08#),
      167 => to_slv(opcode_type, 16#04#),
      168 => to_slv(opcode_type, 16#0D#),
      169 => to_slv(opcode_type, 16#08#),
      170 => to_slv(opcode_type, 16#DE#),
      171 => to_slv(opcode_type, 16#0A#),
      172 => to_slv(opcode_type, 16#09#),
      173 => to_slv(opcode_type, 16#06#),
      174 => to_slv(opcode_type, 16#09#),
      175 => to_slv(opcode_type, 16#10#),
      176 => to_slv(opcode_type, 16#0C#),
      177 => to_slv(opcode_type, 16#07#),
      178 => to_slv(opcode_type, 16#11#),
      179 => to_slv(opcode_type, 16#BA#),
      180 => to_slv(opcode_type, 16#06#),
      181 => to_slv(opcode_type, 16#08#),
      182 => to_slv(opcode_type, 16#0D#),
      183 => to_slv(opcode_type, 16#FD#),
      184 => to_slv(opcode_type, 16#06#),
      185 => to_slv(opcode_type, 16#0E#),
      186 => to_slv(opcode_type, 16#11#),
      187 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#09#),
      193 => to_slv(opcode_type, 16#08#),
      194 => to_slv(opcode_type, 16#04#),
      195 => to_slv(opcode_type, 16#03#),
      196 => to_slv(opcode_type, 16#0E#),
      197 => to_slv(opcode_type, 16#06#),
      198 => to_slv(opcode_type, 16#07#),
      199 => to_slv(opcode_type, 16#0B#),
      200 => to_slv(opcode_type, 16#0C#),
      201 => to_slv(opcode_type, 16#06#),
      202 => to_slv(opcode_type, 16#0E#),
      203 => to_slv(opcode_type, 16#0C#),
      204 => to_slv(opcode_type, 16#07#),
      205 => to_slv(opcode_type, 16#07#),
      206 => to_slv(opcode_type, 16#08#),
      207 => to_slv(opcode_type, 16#0C#),
      208 => to_slv(opcode_type, 16#0E#),
      209 => to_slv(opcode_type, 16#07#),
      210 => to_slv(opcode_type, 16#0E#),
      211 => to_slv(opcode_type, 16#0B#),
      212 => to_slv(opcode_type, 16#08#),
      213 => to_slv(opcode_type, 16#08#),
      214 => to_slv(opcode_type, 16#0D#),
      215 => to_slv(opcode_type, 16#0E#),
      216 => to_slv(opcode_type, 16#09#),
      217 => to_slv(opcode_type, 16#0A#),
      218 => to_slv(opcode_type, 16#48#),
      219 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#08#),
      225 => to_slv(opcode_type, 16#06#),
      226 => to_slv(opcode_type, 16#09#),
      227 => to_slv(opcode_type, 16#05#),
      228 => to_slv(opcode_type, 16#10#),
      229 => to_slv(opcode_type, 16#03#),
      230 => to_slv(opcode_type, 16#0D#),
      231 => to_slv(opcode_type, 16#07#),
      232 => to_slv(opcode_type, 16#04#),
      233 => to_slv(opcode_type, 16#0B#),
      234 => to_slv(opcode_type, 16#05#),
      235 => to_slv(opcode_type, 16#E6#),
      236 => to_slv(opcode_type, 16#09#),
      237 => to_slv(opcode_type, 16#08#),
      238 => to_slv(opcode_type, 16#08#),
      239 => to_slv(opcode_type, 16#0C#),
      240 => to_slv(opcode_type, 16#99#),
      241 => to_slv(opcode_type, 16#07#),
      242 => to_slv(opcode_type, 16#0C#),
      243 => to_slv(opcode_type, 16#0C#),
      244 => to_slv(opcode_type, 16#09#),
      245 => to_slv(opcode_type, 16#06#),
      246 => to_slv(opcode_type, 16#11#),
      247 => to_slv(opcode_type, 16#11#),
      248 => to_slv(opcode_type, 16#08#),
      249 => to_slv(opcode_type, 16#0A#),
      250 => to_slv(opcode_type, 16#0A#),
      251 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#09#),
      257 => to_slv(opcode_type, 16#08#),
      258 => to_slv(opcode_type, 16#02#),
      259 => to_slv(opcode_type, 16#05#),
      260 => to_slv(opcode_type, 16#11#),
      261 => to_slv(opcode_type, 16#07#),
      262 => to_slv(opcode_type, 16#08#),
      263 => to_slv(opcode_type, 16#10#),
      264 => to_slv(opcode_type, 16#7E#),
      265 => to_slv(opcode_type, 16#06#),
      266 => to_slv(opcode_type, 16#0D#),
      267 => to_slv(opcode_type, 16#10#),
      268 => to_slv(opcode_type, 16#08#),
      269 => to_slv(opcode_type, 16#09#),
      270 => to_slv(opcode_type, 16#09#),
      271 => to_slv(opcode_type, 16#8A#),
      272 => to_slv(opcode_type, 16#10#),
      273 => to_slv(opcode_type, 16#06#),
      274 => to_slv(opcode_type, 16#2F#),
      275 => to_slv(opcode_type, 16#0C#),
      276 => to_slv(opcode_type, 16#06#),
      277 => to_slv(opcode_type, 16#06#),
      278 => to_slv(opcode_type, 16#0F#),
      279 => to_slv(opcode_type, 16#10#),
      280 => to_slv(opcode_type, 16#07#),
      281 => to_slv(opcode_type, 16#0D#),
      282 => to_slv(opcode_type, 16#0B#),
      283 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#09#),
      289 => to_slv(opcode_type, 16#08#),
      290 => to_slv(opcode_type, 16#02#),
      291 => to_slv(opcode_type, 16#01#),
      292 => to_slv(opcode_type, 16#0B#),
      293 => to_slv(opcode_type, 16#09#),
      294 => to_slv(opcode_type, 16#07#),
      295 => to_slv(opcode_type, 16#0F#),
      296 => to_slv(opcode_type, 16#99#),
      297 => to_slv(opcode_type, 16#06#),
      298 => to_slv(opcode_type, 16#2B#),
      299 => to_slv(opcode_type, 16#0D#),
      300 => to_slv(opcode_type, 16#06#),
      301 => to_slv(opcode_type, 16#08#),
      302 => to_slv(opcode_type, 16#07#),
      303 => to_slv(opcode_type, 16#0B#),
      304 => to_slv(opcode_type, 16#0B#),
      305 => to_slv(opcode_type, 16#09#),
      306 => to_slv(opcode_type, 16#0C#),
      307 => to_slv(opcode_type, 16#0F#),
      308 => to_slv(opcode_type, 16#06#),
      309 => to_slv(opcode_type, 16#09#),
      310 => to_slv(opcode_type, 16#0E#),
      311 => to_slv(opcode_type, 16#0E#),
      312 => to_slv(opcode_type, 16#06#),
      313 => to_slv(opcode_type, 16#0B#),
      314 => to_slv(opcode_type, 16#0A#),
      315 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#06#),
      321 => to_slv(opcode_type, 16#08#),
      322 => to_slv(opcode_type, 16#02#),
      323 => to_slv(opcode_type, 16#09#),
      324 => to_slv(opcode_type, 16#0F#),
      325 => to_slv(opcode_type, 16#93#),
      326 => to_slv(opcode_type, 16#06#),
      327 => to_slv(opcode_type, 16#08#),
      328 => to_slv(opcode_type, 16#11#),
      329 => to_slv(opcode_type, 16#43#),
      330 => to_slv(opcode_type, 16#07#),
      331 => to_slv(opcode_type, 16#0F#),
      332 => to_slv(opcode_type, 16#2C#),
      333 => to_slv(opcode_type, 16#07#),
      334 => to_slv(opcode_type, 16#08#),
      335 => to_slv(opcode_type, 16#07#),
      336 => to_slv(opcode_type, 16#0A#),
      337 => to_slv(opcode_type, 16#11#),
      338 => to_slv(opcode_type, 16#04#),
      339 => to_slv(opcode_type, 16#10#),
      340 => to_slv(opcode_type, 16#09#),
      341 => to_slv(opcode_type, 16#06#),
      342 => to_slv(opcode_type, 16#0F#),
      343 => to_slv(opcode_type, 16#94#),
      344 => to_slv(opcode_type, 16#09#),
      345 => to_slv(opcode_type, 16#11#),
      346 => to_slv(opcode_type, 16#11#),
      347 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#09#),
      353 => to_slv(opcode_type, 16#06#),
      354 => to_slv(opcode_type, 16#03#),
      355 => to_slv(opcode_type, 16#03#),
      356 => to_slv(opcode_type, 16#0F#),
      357 => to_slv(opcode_type, 16#08#),
      358 => to_slv(opcode_type, 16#07#),
      359 => to_slv(opcode_type, 16#0E#),
      360 => to_slv(opcode_type, 16#0D#),
      361 => to_slv(opcode_type, 16#08#),
      362 => to_slv(opcode_type, 16#11#),
      363 => to_slv(opcode_type, 16#11#),
      364 => to_slv(opcode_type, 16#09#),
      365 => to_slv(opcode_type, 16#06#),
      366 => to_slv(opcode_type, 16#06#),
      367 => to_slv(opcode_type, 16#0E#),
      368 => to_slv(opcode_type, 16#0D#),
      369 => to_slv(opcode_type, 16#07#),
      370 => to_slv(opcode_type, 16#0E#),
      371 => to_slv(opcode_type, 16#0D#),
      372 => to_slv(opcode_type, 16#08#),
      373 => to_slv(opcode_type, 16#07#),
      374 => to_slv(opcode_type, 16#0B#),
      375 => to_slv(opcode_type, 16#0F#),
      376 => to_slv(opcode_type, 16#07#),
      377 => to_slv(opcode_type, 16#11#),
      378 => to_slv(opcode_type, 16#0F#),
      379 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#07#),
      385 => to_slv(opcode_type, 16#07#),
      386 => to_slv(opcode_type, 16#02#),
      387 => to_slv(opcode_type, 16#04#),
      388 => to_slv(opcode_type, 16#0E#),
      389 => to_slv(opcode_type, 16#07#),
      390 => to_slv(opcode_type, 16#09#),
      391 => to_slv(opcode_type, 16#0F#),
      392 => to_slv(opcode_type, 16#42#),
      393 => to_slv(opcode_type, 16#07#),
      394 => to_slv(opcode_type, 16#11#),
      395 => to_slv(opcode_type, 16#10#),
      396 => to_slv(opcode_type, 16#06#),
      397 => to_slv(opcode_type, 16#07#),
      398 => to_slv(opcode_type, 16#06#),
      399 => to_slv(opcode_type, 16#11#),
      400 => to_slv(opcode_type, 16#0D#),
      401 => to_slv(opcode_type, 16#08#),
      402 => to_slv(opcode_type, 16#0B#),
      403 => to_slv(opcode_type, 16#0E#),
      404 => to_slv(opcode_type, 16#06#),
      405 => to_slv(opcode_type, 16#09#),
      406 => to_slv(opcode_type, 16#0C#),
      407 => to_slv(opcode_type, 16#10#),
      408 => to_slv(opcode_type, 16#09#),
      409 => to_slv(opcode_type, 16#11#),
      410 => to_slv(opcode_type, 16#0E#),
      411 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#08#),
      417 => to_slv(opcode_type, 16#06#),
      418 => to_slv(opcode_type, 16#04#),
      419 => to_slv(opcode_type, 16#07#),
      420 => to_slv(opcode_type, 16#0C#),
      421 => to_slv(opcode_type, 16#6A#),
      422 => to_slv(opcode_type, 16#08#),
      423 => to_slv(opcode_type, 16#01#),
      424 => to_slv(opcode_type, 16#0D#),
      425 => to_slv(opcode_type, 16#09#),
      426 => to_slv(opcode_type, 16#0F#),
      427 => to_slv(opcode_type, 16#0F#),
      428 => to_slv(opcode_type, 16#07#),
      429 => to_slv(opcode_type, 16#09#),
      430 => to_slv(opcode_type, 16#07#),
      431 => to_slv(opcode_type, 16#11#),
      432 => to_slv(opcode_type, 16#0B#),
      433 => to_slv(opcode_type, 16#07#),
      434 => to_slv(opcode_type, 16#0B#),
      435 => to_slv(opcode_type, 16#0A#),
      436 => to_slv(opcode_type, 16#08#),
      437 => to_slv(opcode_type, 16#09#),
      438 => to_slv(opcode_type, 16#0C#),
      439 => to_slv(opcode_type, 16#0D#),
      440 => to_slv(opcode_type, 16#09#),
      441 => to_slv(opcode_type, 16#E4#),
      442 => to_slv(opcode_type, 16#0E#),
      443 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#06#),
      449 => to_slv(opcode_type, 16#09#),
      450 => to_slv(opcode_type, 16#09#),
      451 => to_slv(opcode_type, 16#03#),
      452 => to_slv(opcode_type, 16#0F#),
      453 => to_slv(opcode_type, 16#08#),
      454 => to_slv(opcode_type, 16#0E#),
      455 => to_slv(opcode_type, 16#0B#),
      456 => to_slv(opcode_type, 16#02#),
      457 => to_slv(opcode_type, 16#06#),
      458 => to_slv(opcode_type, 16#0E#),
      459 => to_slv(opcode_type, 16#0A#),
      460 => to_slv(opcode_type, 16#07#),
      461 => to_slv(opcode_type, 16#06#),
      462 => to_slv(opcode_type, 16#09#),
      463 => to_slv(opcode_type, 16#0B#),
      464 => to_slv(opcode_type, 16#C8#),
      465 => to_slv(opcode_type, 16#07#),
      466 => to_slv(opcode_type, 16#0C#),
      467 => to_slv(opcode_type, 16#10#),
      468 => to_slv(opcode_type, 16#08#),
      469 => to_slv(opcode_type, 16#08#),
      470 => to_slv(opcode_type, 16#0D#),
      471 => to_slv(opcode_type, 16#0D#),
      472 => to_slv(opcode_type, 16#08#),
      473 => to_slv(opcode_type, 16#10#),
      474 => to_slv(opcode_type, 16#0A#),
      475 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#06#),
      481 => to_slv(opcode_type, 16#07#),
      482 => to_slv(opcode_type, 16#02#),
      483 => to_slv(opcode_type, 16#08#),
      484 => to_slv(opcode_type, 16#0E#),
      485 => to_slv(opcode_type, 16#0E#),
      486 => to_slv(opcode_type, 16#09#),
      487 => to_slv(opcode_type, 16#09#),
      488 => to_slv(opcode_type, 16#10#),
      489 => to_slv(opcode_type, 16#0C#),
      490 => to_slv(opcode_type, 16#02#),
      491 => to_slv(opcode_type, 16#0C#),
      492 => to_slv(opcode_type, 16#07#),
      493 => to_slv(opcode_type, 16#09#),
      494 => to_slv(opcode_type, 16#07#),
      495 => to_slv(opcode_type, 16#0C#),
      496 => to_slv(opcode_type, 16#0E#),
      497 => to_slv(opcode_type, 16#08#),
      498 => to_slv(opcode_type, 16#16#),
      499 => to_slv(opcode_type, 16#2E#),
      500 => to_slv(opcode_type, 16#07#),
      501 => to_slv(opcode_type, 16#07#),
      502 => to_slv(opcode_type, 16#AB#),
      503 => to_slv(opcode_type, 16#0B#),
      504 => to_slv(opcode_type, 16#06#),
      505 => to_slv(opcode_type, 16#47#),
      506 => to_slv(opcode_type, 16#0E#),
      507 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#06#),
      514 => to_slv(opcode_type, 16#03#),
      515 => to_slv(opcode_type, 16#07#),
      516 => to_slv(opcode_type, 16#0E#),
      517 => to_slv(opcode_type, 16#0C#),
      518 => to_slv(opcode_type, 16#06#),
      519 => to_slv(opcode_type, 16#04#),
      520 => to_slv(opcode_type, 16#0A#),
      521 => to_slv(opcode_type, 16#08#),
      522 => to_slv(opcode_type, 16#0C#),
      523 => to_slv(opcode_type, 16#0E#),
      524 => to_slv(opcode_type, 16#08#),
      525 => to_slv(opcode_type, 16#06#),
      526 => to_slv(opcode_type, 16#09#),
      527 => to_slv(opcode_type, 16#0F#),
      528 => to_slv(opcode_type, 16#29#),
      529 => to_slv(opcode_type, 16#08#),
      530 => to_slv(opcode_type, 16#0F#),
      531 => to_slv(opcode_type, 16#10#),
      532 => to_slv(opcode_type, 16#06#),
      533 => to_slv(opcode_type, 16#08#),
      534 => to_slv(opcode_type, 16#10#),
      535 => to_slv(opcode_type, 16#0A#),
      536 => to_slv(opcode_type, 16#06#),
      537 => to_slv(opcode_type, 16#11#),
      538 => to_slv(opcode_type, 16#0E#),
      539 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#09#),
      545 => to_slv(opcode_type, 16#07#),
      546 => to_slv(opcode_type, 16#09#),
      547 => to_slv(opcode_type, 16#01#),
      548 => to_slv(opcode_type, 16#0D#),
      549 => to_slv(opcode_type, 16#07#),
      550 => to_slv(opcode_type, 16#0B#),
      551 => to_slv(opcode_type, 16#0D#),
      552 => to_slv(opcode_type, 16#08#),
      553 => to_slv(opcode_type, 16#07#),
      554 => to_slv(opcode_type, 16#11#),
      555 => to_slv(opcode_type, 16#0D#),
      556 => to_slv(opcode_type, 16#08#),
      557 => to_slv(opcode_type, 16#0D#),
      558 => to_slv(opcode_type, 16#10#),
      559 => to_slv(opcode_type, 16#08#),
      560 => to_slv(opcode_type, 16#04#),
      561 => to_slv(opcode_type, 16#09#),
      562 => to_slv(opcode_type, 16#0D#),
      563 => to_slv(opcode_type, 16#0F#),
      564 => to_slv(opcode_type, 16#08#),
      565 => to_slv(opcode_type, 16#06#),
      566 => to_slv(opcode_type, 16#0F#),
      567 => to_slv(opcode_type, 16#0E#),
      568 => to_slv(opcode_type, 16#07#),
      569 => to_slv(opcode_type, 16#0B#),
      570 => to_slv(opcode_type, 16#0A#),
      571 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#09#),
      577 => to_slv(opcode_type, 16#07#),
      578 => to_slv(opcode_type, 16#04#),
      579 => to_slv(opcode_type, 16#08#),
      580 => to_slv(opcode_type, 16#0A#),
      581 => to_slv(opcode_type, 16#0C#),
      582 => to_slv(opcode_type, 16#07#),
      583 => to_slv(opcode_type, 16#01#),
      584 => to_slv(opcode_type, 16#0D#),
      585 => to_slv(opcode_type, 16#06#),
      586 => to_slv(opcode_type, 16#0F#),
      587 => to_slv(opcode_type, 16#0C#),
      588 => to_slv(opcode_type, 16#09#),
      589 => to_slv(opcode_type, 16#06#),
      590 => to_slv(opcode_type, 16#08#),
      591 => to_slv(opcode_type, 16#0F#),
      592 => to_slv(opcode_type, 16#11#),
      593 => to_slv(opcode_type, 16#06#),
      594 => to_slv(opcode_type, 16#0B#),
      595 => to_slv(opcode_type, 16#0A#),
      596 => to_slv(opcode_type, 16#06#),
      597 => to_slv(opcode_type, 16#08#),
      598 => to_slv(opcode_type, 16#11#),
      599 => to_slv(opcode_type, 16#0D#),
      600 => to_slv(opcode_type, 16#07#),
      601 => to_slv(opcode_type, 16#0A#),
      602 => to_slv(opcode_type, 16#10#),
      603 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#09#),
      609 => to_slv(opcode_type, 16#07#),
      610 => to_slv(opcode_type, 16#03#),
      611 => to_slv(opcode_type, 16#03#),
      612 => to_slv(opcode_type, 16#0A#),
      613 => to_slv(opcode_type, 16#09#),
      614 => to_slv(opcode_type, 16#09#),
      615 => to_slv(opcode_type, 16#0D#),
      616 => to_slv(opcode_type, 16#0B#),
      617 => to_slv(opcode_type, 16#09#),
      618 => to_slv(opcode_type, 16#0E#),
      619 => to_slv(opcode_type, 16#11#),
      620 => to_slv(opcode_type, 16#06#),
      621 => to_slv(opcode_type, 16#09#),
      622 => to_slv(opcode_type, 16#07#),
      623 => to_slv(opcode_type, 16#0E#),
      624 => to_slv(opcode_type, 16#0E#),
      625 => to_slv(opcode_type, 16#07#),
      626 => to_slv(opcode_type, 16#0D#),
      627 => to_slv(opcode_type, 16#8F#),
      628 => to_slv(opcode_type, 16#09#),
      629 => to_slv(opcode_type, 16#07#),
      630 => to_slv(opcode_type, 16#10#),
      631 => to_slv(opcode_type, 16#0D#),
      632 => to_slv(opcode_type, 16#06#),
      633 => to_slv(opcode_type, 16#6D#),
      634 => to_slv(opcode_type, 16#0F#),
      635 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#07#),
      641 => to_slv(opcode_type, 16#08#),
      642 => to_slv(opcode_type, 16#09#),
      643 => to_slv(opcode_type, 16#03#),
      644 => to_slv(opcode_type, 16#0E#),
      645 => to_slv(opcode_type, 16#05#),
      646 => to_slv(opcode_type, 16#FF#),
      647 => to_slv(opcode_type, 16#07#),
      648 => to_slv(opcode_type, 16#04#),
      649 => to_slv(opcode_type, 16#9F#),
      650 => to_slv(opcode_type, 16#08#),
      651 => to_slv(opcode_type, 16#0B#),
      652 => to_slv(opcode_type, 16#0B#),
      653 => to_slv(opcode_type, 16#08#),
      654 => to_slv(opcode_type, 16#07#),
      655 => to_slv(opcode_type, 16#06#),
      656 => to_slv(opcode_type, 16#0C#),
      657 => to_slv(opcode_type, 16#0F#),
      658 => to_slv(opcode_type, 16#03#),
      659 => to_slv(opcode_type, 16#10#),
      660 => to_slv(opcode_type, 16#09#),
      661 => to_slv(opcode_type, 16#08#),
      662 => to_slv(opcode_type, 16#11#),
      663 => to_slv(opcode_type, 16#0D#),
      664 => to_slv(opcode_type, 16#06#),
      665 => to_slv(opcode_type, 16#0E#),
      666 => to_slv(opcode_type, 16#11#),
      667 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#06#),
      673 => to_slv(opcode_type, 16#07#),
      674 => to_slv(opcode_type, 16#09#),
      675 => to_slv(opcode_type, 16#06#),
      676 => to_slv(opcode_type, 16#6C#),
      677 => to_slv(opcode_type, 16#0A#),
      678 => to_slv(opcode_type, 16#03#),
      679 => to_slv(opcode_type, 16#0B#),
      680 => to_slv(opcode_type, 16#01#),
      681 => to_slv(opcode_type, 16#08#),
      682 => to_slv(opcode_type, 16#0B#),
      683 => to_slv(opcode_type, 16#94#),
      684 => to_slv(opcode_type, 16#07#),
      685 => to_slv(opcode_type, 16#08#),
      686 => to_slv(opcode_type, 16#09#),
      687 => to_slv(opcode_type, 16#11#),
      688 => to_slv(opcode_type, 16#0F#),
      689 => to_slv(opcode_type, 16#09#),
      690 => to_slv(opcode_type, 16#0D#),
      691 => to_slv(opcode_type, 16#11#),
      692 => to_slv(opcode_type, 16#09#),
      693 => to_slv(opcode_type, 16#08#),
      694 => to_slv(opcode_type, 16#10#),
      695 => to_slv(opcode_type, 16#0D#),
      696 => to_slv(opcode_type, 16#09#),
      697 => to_slv(opcode_type, 16#11#),
      698 => to_slv(opcode_type, 16#0C#),
      699 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#08#),
      705 => to_slv(opcode_type, 16#08#),
      706 => to_slv(opcode_type, 16#04#),
      707 => to_slv(opcode_type, 16#09#),
      708 => to_slv(opcode_type, 16#0B#),
      709 => to_slv(opcode_type, 16#0B#),
      710 => to_slv(opcode_type, 16#09#),
      711 => to_slv(opcode_type, 16#01#),
      712 => to_slv(opcode_type, 16#0A#),
      713 => to_slv(opcode_type, 16#09#),
      714 => to_slv(opcode_type, 16#0C#),
      715 => to_slv(opcode_type, 16#0A#),
      716 => to_slv(opcode_type, 16#07#),
      717 => to_slv(opcode_type, 16#06#),
      718 => to_slv(opcode_type, 16#09#),
      719 => to_slv(opcode_type, 16#0B#),
      720 => to_slv(opcode_type, 16#0A#),
      721 => to_slv(opcode_type, 16#09#),
      722 => to_slv(opcode_type, 16#0B#),
      723 => to_slv(opcode_type, 16#0E#),
      724 => to_slv(opcode_type, 16#08#),
      725 => to_slv(opcode_type, 16#08#),
      726 => to_slv(opcode_type, 16#0A#),
      727 => to_slv(opcode_type, 16#0A#),
      728 => to_slv(opcode_type, 16#06#),
      729 => to_slv(opcode_type, 16#0C#),
      730 => to_slv(opcode_type, 16#0B#),
      731 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#08#),
      737 => to_slv(opcode_type, 16#09#),
      738 => to_slv(opcode_type, 16#09#),
      739 => to_slv(opcode_type, 16#07#),
      740 => to_slv(opcode_type, 16#11#),
      741 => to_slv(opcode_type, 16#11#),
      742 => to_slv(opcode_type, 16#04#),
      743 => to_slv(opcode_type, 16#0E#),
      744 => to_slv(opcode_type, 16#02#),
      745 => to_slv(opcode_type, 16#09#),
      746 => to_slv(opcode_type, 16#91#),
      747 => to_slv(opcode_type, 16#0D#),
      748 => to_slv(opcode_type, 16#09#),
      749 => to_slv(opcode_type, 16#08#),
      750 => to_slv(opcode_type, 16#09#),
      751 => to_slv(opcode_type, 16#0D#),
      752 => to_slv(opcode_type, 16#11#),
      753 => to_slv(opcode_type, 16#06#),
      754 => to_slv(opcode_type, 16#0A#),
      755 => to_slv(opcode_type, 16#0F#),
      756 => to_slv(opcode_type, 16#09#),
      757 => to_slv(opcode_type, 16#08#),
      758 => to_slv(opcode_type, 16#0B#),
      759 => to_slv(opcode_type, 16#0C#),
      760 => to_slv(opcode_type, 16#06#),
      761 => to_slv(opcode_type, 16#77#),
      762 => to_slv(opcode_type, 16#10#),
      763 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#08#),
      769 => to_slv(opcode_type, 16#09#),
      770 => to_slv(opcode_type, 16#07#),
      771 => to_slv(opcode_type, 16#07#),
      772 => to_slv(opcode_type, 16#0B#),
      773 => to_slv(opcode_type, 16#11#),
      774 => to_slv(opcode_type, 16#01#),
      775 => to_slv(opcode_type, 16#0E#),
      776 => to_slv(opcode_type, 16#04#),
      777 => to_slv(opcode_type, 16#07#),
      778 => to_slv(opcode_type, 16#0B#),
      779 => to_slv(opcode_type, 16#0A#),
      780 => to_slv(opcode_type, 16#08#),
      781 => to_slv(opcode_type, 16#08#),
      782 => to_slv(opcode_type, 16#09#),
      783 => to_slv(opcode_type, 16#0C#),
      784 => to_slv(opcode_type, 16#0C#),
      785 => to_slv(opcode_type, 16#08#),
      786 => to_slv(opcode_type, 16#0E#),
      787 => to_slv(opcode_type, 16#0D#),
      788 => to_slv(opcode_type, 16#09#),
      789 => to_slv(opcode_type, 16#08#),
      790 => to_slv(opcode_type, 16#0F#),
      791 => to_slv(opcode_type, 16#0E#),
      792 => to_slv(opcode_type, 16#07#),
      793 => to_slv(opcode_type, 16#0B#),
      794 => to_slv(opcode_type, 16#11#),
      795 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#07#),
      801 => to_slv(opcode_type, 16#06#),
      802 => to_slv(opcode_type, 16#03#),
      803 => to_slv(opcode_type, 16#09#),
      804 => to_slv(opcode_type, 16#10#),
      805 => to_slv(opcode_type, 16#E4#),
      806 => to_slv(opcode_type, 16#09#),
      807 => to_slv(opcode_type, 16#02#),
      808 => to_slv(opcode_type, 16#0A#),
      809 => to_slv(opcode_type, 16#07#),
      810 => to_slv(opcode_type, 16#0A#),
      811 => to_slv(opcode_type, 16#0B#),
      812 => to_slv(opcode_type, 16#07#),
      813 => to_slv(opcode_type, 16#08#),
      814 => to_slv(opcode_type, 16#07#),
      815 => to_slv(opcode_type, 16#10#),
      816 => to_slv(opcode_type, 16#11#),
      817 => to_slv(opcode_type, 16#08#),
      818 => to_slv(opcode_type, 16#77#),
      819 => to_slv(opcode_type, 16#0A#),
      820 => to_slv(opcode_type, 16#06#),
      821 => to_slv(opcode_type, 16#06#),
      822 => to_slv(opcode_type, 16#8C#),
      823 => to_slv(opcode_type, 16#11#),
      824 => to_slv(opcode_type, 16#06#),
      825 => to_slv(opcode_type, 16#0F#),
      826 => to_slv(opcode_type, 16#0F#),
      827 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#06#),
      833 => to_slv(opcode_type, 16#09#),
      834 => to_slv(opcode_type, 16#02#),
      835 => to_slv(opcode_type, 16#03#),
      836 => to_slv(opcode_type, 16#10#),
      837 => to_slv(opcode_type, 16#06#),
      838 => to_slv(opcode_type, 16#08#),
      839 => to_slv(opcode_type, 16#0F#),
      840 => to_slv(opcode_type, 16#10#),
      841 => to_slv(opcode_type, 16#09#),
      842 => to_slv(opcode_type, 16#0A#),
      843 => to_slv(opcode_type, 16#11#),
      844 => to_slv(opcode_type, 16#07#),
      845 => to_slv(opcode_type, 16#09#),
      846 => to_slv(opcode_type, 16#06#),
      847 => to_slv(opcode_type, 16#0C#),
      848 => to_slv(opcode_type, 16#10#),
      849 => to_slv(opcode_type, 16#08#),
      850 => to_slv(opcode_type, 16#0B#),
      851 => to_slv(opcode_type, 16#10#),
      852 => to_slv(opcode_type, 16#07#),
      853 => to_slv(opcode_type, 16#07#),
      854 => to_slv(opcode_type, 16#0E#),
      855 => to_slv(opcode_type, 16#0D#),
      856 => to_slv(opcode_type, 16#07#),
      857 => to_slv(opcode_type, 16#47#),
      858 => to_slv(opcode_type, 16#10#),
      859 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#07#),
      865 => to_slv(opcode_type, 16#09#),
      866 => to_slv(opcode_type, 16#05#),
      867 => to_slv(opcode_type, 16#02#),
      868 => to_slv(opcode_type, 16#0A#),
      869 => to_slv(opcode_type, 16#09#),
      870 => to_slv(opcode_type, 16#08#),
      871 => to_slv(opcode_type, 16#0E#),
      872 => to_slv(opcode_type, 16#0F#),
      873 => to_slv(opcode_type, 16#08#),
      874 => to_slv(opcode_type, 16#0A#),
      875 => to_slv(opcode_type, 16#0D#),
      876 => to_slv(opcode_type, 16#08#),
      877 => to_slv(opcode_type, 16#08#),
      878 => to_slv(opcode_type, 16#07#),
      879 => to_slv(opcode_type, 16#0A#),
      880 => to_slv(opcode_type, 16#11#),
      881 => to_slv(opcode_type, 16#09#),
      882 => to_slv(opcode_type, 16#0A#),
      883 => to_slv(opcode_type, 16#0C#),
      884 => to_slv(opcode_type, 16#06#),
      885 => to_slv(opcode_type, 16#08#),
      886 => to_slv(opcode_type, 16#0E#),
      887 => to_slv(opcode_type, 16#10#),
      888 => to_slv(opcode_type, 16#09#),
      889 => to_slv(opcode_type, 16#A4#),
      890 => to_slv(opcode_type, 16#0F#),
      891 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#08#),
      897 => to_slv(opcode_type, 16#09#),
      898 => to_slv(opcode_type, 16#09#),
      899 => to_slv(opcode_type, 16#06#),
      900 => to_slv(opcode_type, 16#0B#),
      901 => to_slv(opcode_type, 16#0B#),
      902 => to_slv(opcode_type, 16#02#),
      903 => to_slv(opcode_type, 16#0C#),
      904 => to_slv(opcode_type, 16#06#),
      905 => to_slv(opcode_type, 16#02#),
      906 => to_slv(opcode_type, 16#0F#),
      907 => to_slv(opcode_type, 16#06#),
      908 => to_slv(opcode_type, 16#0B#),
      909 => to_slv(opcode_type, 16#0C#),
      910 => to_slv(opcode_type, 16#07#),
      911 => to_slv(opcode_type, 16#09#),
      912 => to_slv(opcode_type, 16#06#),
      913 => to_slv(opcode_type, 16#0A#),
      914 => to_slv(opcode_type, 16#0C#),
      915 => to_slv(opcode_type, 16#06#),
      916 => to_slv(opcode_type, 16#11#),
      917 => to_slv(opcode_type, 16#0B#),
      918 => to_slv(opcode_type, 16#06#),
      919 => to_slv(opcode_type, 16#09#),
      920 => to_slv(opcode_type, 16#11#),
      921 => to_slv(opcode_type, 16#10#),
      922 => to_slv(opcode_type, 16#11#),
      923 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#09#),
      929 => to_slv(opcode_type, 16#07#),
      930 => to_slv(opcode_type, 16#06#),
      931 => to_slv(opcode_type, 16#01#),
      932 => to_slv(opcode_type, 16#0B#),
      933 => to_slv(opcode_type, 16#04#),
      934 => to_slv(opcode_type, 16#0B#),
      935 => to_slv(opcode_type, 16#07#),
      936 => to_slv(opcode_type, 16#04#),
      937 => to_slv(opcode_type, 16#0E#),
      938 => to_slv(opcode_type, 16#05#),
      939 => to_slv(opcode_type, 16#0A#),
      940 => to_slv(opcode_type, 16#07#),
      941 => to_slv(opcode_type, 16#06#),
      942 => to_slv(opcode_type, 16#08#),
      943 => to_slv(opcode_type, 16#0D#),
      944 => to_slv(opcode_type, 16#0D#),
      945 => to_slv(opcode_type, 16#08#),
      946 => to_slv(opcode_type, 16#10#),
      947 => to_slv(opcode_type, 16#0D#),
      948 => to_slv(opcode_type, 16#07#),
      949 => to_slv(opcode_type, 16#07#),
      950 => to_slv(opcode_type, 16#6F#),
      951 => to_slv(opcode_type, 16#0C#),
      952 => to_slv(opcode_type, 16#07#),
      953 => to_slv(opcode_type, 16#10#),
      954 => to_slv(opcode_type, 16#0C#),
      955 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#07#),
      962 => to_slv(opcode_type, 16#03#),
      963 => to_slv(opcode_type, 16#01#),
      964 => to_slv(opcode_type, 16#0E#),
      965 => to_slv(opcode_type, 16#09#),
      966 => to_slv(opcode_type, 16#08#),
      967 => to_slv(opcode_type, 16#0D#),
      968 => to_slv(opcode_type, 16#0E#),
      969 => to_slv(opcode_type, 16#09#),
      970 => to_slv(opcode_type, 16#10#),
      971 => to_slv(opcode_type, 16#FD#),
      972 => to_slv(opcode_type, 16#06#),
      973 => to_slv(opcode_type, 16#07#),
      974 => to_slv(opcode_type, 16#08#),
      975 => to_slv(opcode_type, 16#0F#),
      976 => to_slv(opcode_type, 16#0A#),
      977 => to_slv(opcode_type, 16#06#),
      978 => to_slv(opcode_type, 16#0B#),
      979 => to_slv(opcode_type, 16#11#),
      980 => to_slv(opcode_type, 16#09#),
      981 => to_slv(opcode_type, 16#06#),
      982 => to_slv(opcode_type, 16#0A#),
      983 => to_slv(opcode_type, 16#11#),
      984 => to_slv(opcode_type, 16#08#),
      985 => to_slv(opcode_type, 16#0D#),
      986 => to_slv(opcode_type, 16#0E#),
      987 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#09#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#05#),
      995 => to_slv(opcode_type, 16#02#),
      996 => to_slv(opcode_type, 16#0D#),
      997 => to_slv(opcode_type, 16#07#),
      998 => to_slv(opcode_type, 16#08#),
      999 => to_slv(opcode_type, 16#0A#),
      1000 => to_slv(opcode_type, 16#0F#),
      1001 => to_slv(opcode_type, 16#09#),
      1002 => to_slv(opcode_type, 16#0A#),
      1003 => to_slv(opcode_type, 16#0F#),
      1004 => to_slv(opcode_type, 16#06#),
      1005 => to_slv(opcode_type, 16#08#),
      1006 => to_slv(opcode_type, 16#09#),
      1007 => to_slv(opcode_type, 16#0F#),
      1008 => to_slv(opcode_type, 16#0C#),
      1009 => to_slv(opcode_type, 16#07#),
      1010 => to_slv(opcode_type, 16#0E#),
      1011 => to_slv(opcode_type, 16#10#),
      1012 => to_slv(opcode_type, 16#08#),
      1013 => to_slv(opcode_type, 16#09#),
      1014 => to_slv(opcode_type, 16#0D#),
      1015 => to_slv(opcode_type, 16#0C#),
      1016 => to_slv(opcode_type, 16#06#),
      1017 => to_slv(opcode_type, 16#0F#),
      1018 => to_slv(opcode_type, 16#10#),
      1019 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#08#),
      1025 => to_slv(opcode_type, 16#08#),
      1026 => to_slv(opcode_type, 16#07#),
      1027 => to_slv(opcode_type, 16#08#),
      1028 => to_slv(opcode_type, 16#9B#),
      1029 => to_slv(opcode_type, 16#0C#),
      1030 => to_slv(opcode_type, 16#01#),
      1031 => to_slv(opcode_type, 16#10#),
      1032 => to_slv(opcode_type, 16#03#),
      1033 => to_slv(opcode_type, 16#07#),
      1034 => to_slv(opcode_type, 16#0A#),
      1035 => to_slv(opcode_type, 16#97#),
      1036 => to_slv(opcode_type, 16#09#),
      1037 => to_slv(opcode_type, 16#06#),
      1038 => to_slv(opcode_type, 16#07#),
      1039 => to_slv(opcode_type, 16#10#),
      1040 => to_slv(opcode_type, 16#10#),
      1041 => to_slv(opcode_type, 16#09#),
      1042 => to_slv(opcode_type, 16#0F#),
      1043 => to_slv(opcode_type, 16#0E#),
      1044 => to_slv(opcode_type, 16#09#),
      1045 => to_slv(opcode_type, 16#09#),
      1046 => to_slv(opcode_type, 16#10#),
      1047 => to_slv(opcode_type, 16#0A#),
      1048 => to_slv(opcode_type, 16#06#),
      1049 => to_slv(opcode_type, 16#0B#),
      1050 => to_slv(opcode_type, 16#10#),
      1051 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#06#),
      1057 => to_slv(opcode_type, 16#06#),
      1058 => to_slv(opcode_type, 16#07#),
      1059 => to_slv(opcode_type, 16#01#),
      1060 => to_slv(opcode_type, 16#0E#),
      1061 => to_slv(opcode_type, 16#01#),
      1062 => to_slv(opcode_type, 16#10#),
      1063 => to_slv(opcode_type, 16#06#),
      1064 => to_slv(opcode_type, 16#01#),
      1065 => to_slv(opcode_type, 16#0A#),
      1066 => to_slv(opcode_type, 16#06#),
      1067 => to_slv(opcode_type, 16#0B#),
      1068 => to_slv(opcode_type, 16#0B#),
      1069 => to_slv(opcode_type, 16#06#),
      1070 => to_slv(opcode_type, 16#09#),
      1071 => to_slv(opcode_type, 16#04#),
      1072 => to_slv(opcode_type, 16#0C#),
      1073 => to_slv(opcode_type, 16#08#),
      1074 => to_slv(opcode_type, 16#AA#),
      1075 => to_slv(opcode_type, 16#0F#),
      1076 => to_slv(opcode_type, 16#09#),
      1077 => to_slv(opcode_type, 16#08#),
      1078 => to_slv(opcode_type, 16#10#),
      1079 => to_slv(opcode_type, 16#10#),
      1080 => to_slv(opcode_type, 16#08#),
      1081 => to_slv(opcode_type, 16#0F#),
      1082 => to_slv(opcode_type, 16#AC#),
      1083 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#09#),
      1089 => to_slv(opcode_type, 16#08#),
      1090 => to_slv(opcode_type, 16#09#),
      1091 => to_slv(opcode_type, 16#07#),
      1092 => to_slv(opcode_type, 16#0B#),
      1093 => to_slv(opcode_type, 16#0C#),
      1094 => to_slv(opcode_type, 16#02#),
      1095 => to_slv(opcode_type, 16#0C#),
      1096 => to_slv(opcode_type, 16#05#),
      1097 => to_slv(opcode_type, 16#06#),
      1098 => to_slv(opcode_type, 16#10#),
      1099 => to_slv(opcode_type, 16#10#),
      1100 => to_slv(opcode_type, 16#09#),
      1101 => to_slv(opcode_type, 16#07#),
      1102 => to_slv(opcode_type, 16#09#),
      1103 => to_slv(opcode_type, 16#10#),
      1104 => to_slv(opcode_type, 16#0E#),
      1105 => to_slv(opcode_type, 16#08#),
      1106 => to_slv(opcode_type, 16#11#),
      1107 => to_slv(opcode_type, 16#11#),
      1108 => to_slv(opcode_type, 16#09#),
      1109 => to_slv(opcode_type, 16#08#),
      1110 => to_slv(opcode_type, 16#0B#),
      1111 => to_slv(opcode_type, 16#0D#),
      1112 => to_slv(opcode_type, 16#09#),
      1113 => to_slv(opcode_type, 16#0E#),
      1114 => to_slv(opcode_type, 16#0D#),
      1115 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#08#),
      1121 => to_slv(opcode_type, 16#08#),
      1122 => to_slv(opcode_type, 16#04#),
      1123 => to_slv(opcode_type, 16#06#),
      1124 => to_slv(opcode_type, 16#0A#),
      1125 => to_slv(opcode_type, 16#0A#),
      1126 => to_slv(opcode_type, 16#06#),
      1127 => to_slv(opcode_type, 16#09#),
      1128 => to_slv(opcode_type, 16#11#),
      1129 => to_slv(opcode_type, 16#0E#),
      1130 => to_slv(opcode_type, 16#08#),
      1131 => to_slv(opcode_type, 16#0B#),
      1132 => to_slv(opcode_type, 16#10#),
      1133 => to_slv(opcode_type, 16#08#),
      1134 => to_slv(opcode_type, 16#09#),
      1135 => to_slv(opcode_type, 16#02#),
      1136 => to_slv(opcode_type, 16#11#),
      1137 => to_slv(opcode_type, 16#08#),
      1138 => to_slv(opcode_type, 16#0C#),
      1139 => to_slv(opcode_type, 16#0C#),
      1140 => to_slv(opcode_type, 16#09#),
      1141 => to_slv(opcode_type, 16#06#),
      1142 => to_slv(opcode_type, 16#0F#),
      1143 => to_slv(opcode_type, 16#4F#),
      1144 => to_slv(opcode_type, 16#06#),
      1145 => to_slv(opcode_type, 16#E4#),
      1146 => to_slv(opcode_type, 16#0D#),
      1147 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#08#),
      1153 => to_slv(opcode_type, 16#06#),
      1154 => to_slv(opcode_type, 16#04#),
      1155 => to_slv(opcode_type, 16#04#),
      1156 => to_slv(opcode_type, 16#0B#),
      1157 => to_slv(opcode_type, 16#07#),
      1158 => to_slv(opcode_type, 16#08#),
      1159 => to_slv(opcode_type, 16#91#),
      1160 => to_slv(opcode_type, 16#0B#),
      1161 => to_slv(opcode_type, 16#06#),
      1162 => to_slv(opcode_type, 16#0B#),
      1163 => to_slv(opcode_type, 16#11#),
      1164 => to_slv(opcode_type, 16#07#),
      1165 => to_slv(opcode_type, 16#06#),
      1166 => to_slv(opcode_type, 16#06#),
      1167 => to_slv(opcode_type, 16#0B#),
      1168 => to_slv(opcode_type, 16#0B#),
      1169 => to_slv(opcode_type, 16#06#),
      1170 => to_slv(opcode_type, 16#0D#),
      1171 => to_slv(opcode_type, 16#11#),
      1172 => to_slv(opcode_type, 16#09#),
      1173 => to_slv(opcode_type, 16#06#),
      1174 => to_slv(opcode_type, 16#0B#),
      1175 => to_slv(opcode_type, 16#FA#),
      1176 => to_slv(opcode_type, 16#07#),
      1177 => to_slv(opcode_type, 16#10#),
      1178 => to_slv(opcode_type, 16#10#),
      1179 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#06#),
      1185 => to_slv(opcode_type, 16#08#),
      1186 => to_slv(opcode_type, 16#04#),
      1187 => to_slv(opcode_type, 16#05#),
      1188 => to_slv(opcode_type, 16#10#),
      1189 => to_slv(opcode_type, 16#09#),
      1190 => to_slv(opcode_type, 16#07#),
      1191 => to_slv(opcode_type, 16#0D#),
      1192 => to_slv(opcode_type, 16#0C#),
      1193 => to_slv(opcode_type, 16#09#),
      1194 => to_slv(opcode_type, 16#0E#),
      1195 => to_slv(opcode_type, 16#0F#),
      1196 => to_slv(opcode_type, 16#07#),
      1197 => to_slv(opcode_type, 16#09#),
      1198 => to_slv(opcode_type, 16#06#),
      1199 => to_slv(opcode_type, 16#48#),
      1200 => to_slv(opcode_type, 16#0E#),
      1201 => to_slv(opcode_type, 16#09#),
      1202 => to_slv(opcode_type, 16#11#),
      1203 => to_slv(opcode_type, 16#0E#),
      1204 => to_slv(opcode_type, 16#08#),
      1205 => to_slv(opcode_type, 16#07#),
      1206 => to_slv(opcode_type, 16#0B#),
      1207 => to_slv(opcode_type, 16#11#),
      1208 => to_slv(opcode_type, 16#08#),
      1209 => to_slv(opcode_type, 16#BC#),
      1210 => to_slv(opcode_type, 16#0D#),
      1211 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#09#),
      1217 => to_slv(opcode_type, 16#08#),
      1218 => to_slv(opcode_type, 16#09#),
      1219 => to_slv(opcode_type, 16#09#),
      1220 => to_slv(opcode_type, 16#11#),
      1221 => to_slv(opcode_type, 16#0F#),
      1222 => to_slv(opcode_type, 16#03#),
      1223 => to_slv(opcode_type, 16#0F#),
      1224 => to_slv(opcode_type, 16#05#),
      1225 => to_slv(opcode_type, 16#08#),
      1226 => to_slv(opcode_type, 16#0B#),
      1227 => to_slv(opcode_type, 16#0C#),
      1228 => to_slv(opcode_type, 16#07#),
      1229 => to_slv(opcode_type, 16#06#),
      1230 => to_slv(opcode_type, 16#07#),
      1231 => to_slv(opcode_type, 16#10#),
      1232 => to_slv(opcode_type, 16#0B#),
      1233 => to_slv(opcode_type, 16#06#),
      1234 => to_slv(opcode_type, 16#37#),
      1235 => to_slv(opcode_type, 16#0B#),
      1236 => to_slv(opcode_type, 16#06#),
      1237 => to_slv(opcode_type, 16#09#),
      1238 => to_slv(opcode_type, 16#0E#),
      1239 => to_slv(opcode_type, 16#0C#),
      1240 => to_slv(opcode_type, 16#06#),
      1241 => to_slv(opcode_type, 16#0F#),
      1242 => to_slv(opcode_type, 16#11#),
      1243 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#07#),
      1249 => to_slv(opcode_type, 16#09#),
      1250 => to_slv(opcode_type, 16#09#),
      1251 => to_slv(opcode_type, 16#09#),
      1252 => to_slv(opcode_type, 16#0D#),
      1253 => to_slv(opcode_type, 16#0B#),
      1254 => to_slv(opcode_type, 16#09#),
      1255 => to_slv(opcode_type, 16#B6#),
      1256 => to_slv(opcode_type, 16#0E#),
      1257 => to_slv(opcode_type, 16#03#),
      1258 => to_slv(opcode_type, 16#08#),
      1259 => to_slv(opcode_type, 16#0A#),
      1260 => to_slv(opcode_type, 16#0B#),
      1261 => to_slv(opcode_type, 16#07#),
      1262 => to_slv(opcode_type, 16#06#),
      1263 => to_slv(opcode_type, 16#02#),
      1264 => to_slv(opcode_type, 16#0F#),
      1265 => to_slv(opcode_type, 16#09#),
      1266 => to_slv(opcode_type, 16#0C#),
      1267 => to_slv(opcode_type, 16#0F#),
      1268 => to_slv(opcode_type, 16#07#),
      1269 => to_slv(opcode_type, 16#09#),
      1270 => to_slv(opcode_type, 16#11#),
      1271 => to_slv(opcode_type, 16#0F#),
      1272 => to_slv(opcode_type, 16#09#),
      1273 => to_slv(opcode_type, 16#50#),
      1274 => to_slv(opcode_type, 16#0B#),
      1275 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#09#),
      1282 => to_slv(opcode_type, 16#08#),
      1283 => to_slv(opcode_type, 16#05#),
      1284 => to_slv(opcode_type, 16#0C#),
      1285 => to_slv(opcode_type, 16#09#),
      1286 => to_slv(opcode_type, 16#0F#),
      1287 => to_slv(opcode_type, 16#10#),
      1288 => to_slv(opcode_type, 16#07#),
      1289 => to_slv(opcode_type, 16#06#),
      1290 => to_slv(opcode_type, 16#14#),
      1291 => to_slv(opcode_type, 16#10#),
      1292 => to_slv(opcode_type, 16#06#),
      1293 => to_slv(opcode_type, 16#0C#),
      1294 => to_slv(opcode_type, 16#0B#),
      1295 => to_slv(opcode_type, 16#07#),
      1296 => to_slv(opcode_type, 16#08#),
      1297 => to_slv(opcode_type, 16#02#),
      1298 => to_slv(opcode_type, 16#10#),
      1299 => to_slv(opcode_type, 16#03#),
      1300 => to_slv(opcode_type, 16#0C#),
      1301 => to_slv(opcode_type, 16#06#),
      1302 => to_slv(opcode_type, 16#03#),
      1303 => to_slv(opcode_type, 16#10#),
      1304 => to_slv(opcode_type, 16#07#),
      1305 => to_slv(opcode_type, 16#0B#),
      1306 => to_slv(opcode_type, 16#11#),
      1307 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#09#),
      1313 => to_slv(opcode_type, 16#08#),
      1314 => to_slv(opcode_type, 16#05#),
      1315 => to_slv(opcode_type, 16#08#),
      1316 => to_slv(opcode_type, 16#11#),
      1317 => to_slv(opcode_type, 16#0D#),
      1318 => to_slv(opcode_type, 16#08#),
      1319 => to_slv(opcode_type, 16#02#),
      1320 => to_slv(opcode_type, 16#0F#),
      1321 => to_slv(opcode_type, 16#07#),
      1322 => to_slv(opcode_type, 16#0A#),
      1323 => to_slv(opcode_type, 16#11#),
      1324 => to_slv(opcode_type, 16#06#),
      1325 => to_slv(opcode_type, 16#06#),
      1326 => to_slv(opcode_type, 16#09#),
      1327 => to_slv(opcode_type, 16#0F#),
      1328 => to_slv(opcode_type, 16#0C#),
      1329 => to_slv(opcode_type, 16#08#),
      1330 => to_slv(opcode_type, 16#0F#),
      1331 => to_slv(opcode_type, 16#0F#),
      1332 => to_slv(opcode_type, 16#07#),
      1333 => to_slv(opcode_type, 16#06#),
      1334 => to_slv(opcode_type, 16#10#),
      1335 => to_slv(opcode_type, 16#10#),
      1336 => to_slv(opcode_type, 16#09#),
      1337 => to_slv(opcode_type, 16#0F#),
      1338 => to_slv(opcode_type, 16#10#),
      1339 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#06#),
      1345 => to_slv(opcode_type, 16#06#),
      1346 => to_slv(opcode_type, 16#08#),
      1347 => to_slv(opcode_type, 16#02#),
      1348 => to_slv(opcode_type, 16#0B#),
      1349 => to_slv(opcode_type, 16#08#),
      1350 => to_slv(opcode_type, 16#90#),
      1351 => to_slv(opcode_type, 16#0F#),
      1352 => to_slv(opcode_type, 16#08#),
      1353 => to_slv(opcode_type, 16#09#),
      1354 => to_slv(opcode_type, 16#0B#),
      1355 => to_slv(opcode_type, 16#11#),
      1356 => to_slv(opcode_type, 16#05#),
      1357 => to_slv(opcode_type, 16#0E#),
      1358 => to_slv(opcode_type, 16#08#),
      1359 => to_slv(opcode_type, 16#08#),
      1360 => to_slv(opcode_type, 16#04#),
      1361 => to_slv(opcode_type, 16#10#),
      1362 => to_slv(opcode_type, 16#04#),
      1363 => to_slv(opcode_type, 16#83#),
      1364 => to_slv(opcode_type, 16#06#),
      1365 => to_slv(opcode_type, 16#08#),
      1366 => to_slv(opcode_type, 16#0F#),
      1367 => to_slv(opcode_type, 16#0D#),
      1368 => to_slv(opcode_type, 16#09#),
      1369 => to_slv(opcode_type, 16#22#),
      1370 => to_slv(opcode_type, 16#0A#),
      1371 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#07#),
      1377 => to_slv(opcode_type, 16#07#),
      1378 => to_slv(opcode_type, 16#01#),
      1379 => to_slv(opcode_type, 16#02#),
      1380 => to_slv(opcode_type, 16#0F#),
      1381 => to_slv(opcode_type, 16#06#),
      1382 => to_slv(opcode_type, 16#07#),
      1383 => to_slv(opcode_type, 16#11#),
      1384 => to_slv(opcode_type, 16#11#),
      1385 => to_slv(opcode_type, 16#09#),
      1386 => to_slv(opcode_type, 16#0C#),
      1387 => to_slv(opcode_type, 16#10#),
      1388 => to_slv(opcode_type, 16#07#),
      1389 => to_slv(opcode_type, 16#09#),
      1390 => to_slv(opcode_type, 16#06#),
      1391 => to_slv(opcode_type, 16#0C#),
      1392 => to_slv(opcode_type, 16#0F#),
      1393 => to_slv(opcode_type, 16#09#),
      1394 => to_slv(opcode_type, 16#11#),
      1395 => to_slv(opcode_type, 16#0D#),
      1396 => to_slv(opcode_type, 16#09#),
      1397 => to_slv(opcode_type, 16#06#),
      1398 => to_slv(opcode_type, 16#11#),
      1399 => to_slv(opcode_type, 16#0E#),
      1400 => to_slv(opcode_type, 16#06#),
      1401 => to_slv(opcode_type, 16#0D#),
      1402 => to_slv(opcode_type, 16#0D#),
      1403 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#07#),
      1409 => to_slv(opcode_type, 16#07#),
      1410 => to_slv(opcode_type, 16#07#),
      1411 => to_slv(opcode_type, 16#06#),
      1412 => to_slv(opcode_type, 16#0F#),
      1413 => to_slv(opcode_type, 16#0A#),
      1414 => to_slv(opcode_type, 16#06#),
      1415 => to_slv(opcode_type, 16#0B#),
      1416 => to_slv(opcode_type, 16#0D#),
      1417 => to_slv(opcode_type, 16#01#),
      1418 => to_slv(opcode_type, 16#04#),
      1419 => to_slv(opcode_type, 16#0A#),
      1420 => to_slv(opcode_type, 16#07#),
      1421 => to_slv(opcode_type, 16#09#),
      1422 => to_slv(opcode_type, 16#06#),
      1423 => to_slv(opcode_type, 16#10#),
      1424 => to_slv(opcode_type, 16#0E#),
      1425 => to_slv(opcode_type, 16#09#),
      1426 => to_slv(opcode_type, 16#11#),
      1427 => to_slv(opcode_type, 16#0A#),
      1428 => to_slv(opcode_type, 16#06#),
      1429 => to_slv(opcode_type, 16#08#),
      1430 => to_slv(opcode_type, 16#11#),
      1431 => to_slv(opcode_type, 16#10#),
      1432 => to_slv(opcode_type, 16#07#),
      1433 => to_slv(opcode_type, 16#0E#),
      1434 => to_slv(opcode_type, 16#11#),
      1435 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#06#),
      1441 => to_slv(opcode_type, 16#09#),
      1442 => to_slv(opcode_type, 16#03#),
      1443 => to_slv(opcode_type, 16#09#),
      1444 => to_slv(opcode_type, 16#10#),
      1445 => to_slv(opcode_type, 16#0D#),
      1446 => to_slv(opcode_type, 16#08#),
      1447 => to_slv(opcode_type, 16#06#),
      1448 => to_slv(opcode_type, 16#0F#),
      1449 => to_slv(opcode_type, 16#61#),
      1450 => to_slv(opcode_type, 16#09#),
      1451 => to_slv(opcode_type, 16#0C#),
      1452 => to_slv(opcode_type, 16#0C#),
      1453 => to_slv(opcode_type, 16#06#),
      1454 => to_slv(opcode_type, 16#09#),
      1455 => to_slv(opcode_type, 16#04#),
      1456 => to_slv(opcode_type, 16#11#),
      1457 => to_slv(opcode_type, 16#06#),
      1458 => to_slv(opcode_type, 16#A6#),
      1459 => to_slv(opcode_type, 16#0A#),
      1460 => to_slv(opcode_type, 16#06#),
      1461 => to_slv(opcode_type, 16#07#),
      1462 => to_slv(opcode_type, 16#0F#),
      1463 => to_slv(opcode_type, 16#0B#),
      1464 => to_slv(opcode_type, 16#09#),
      1465 => to_slv(opcode_type, 16#0F#),
      1466 => to_slv(opcode_type, 16#11#),
      1467 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#06#),
      1473 => to_slv(opcode_type, 16#07#),
      1474 => to_slv(opcode_type, 16#05#),
      1475 => to_slv(opcode_type, 16#09#),
      1476 => to_slv(opcode_type, 16#0C#),
      1477 => to_slv(opcode_type, 16#0A#),
      1478 => to_slv(opcode_type, 16#08#),
      1479 => to_slv(opcode_type, 16#08#),
      1480 => to_slv(opcode_type, 16#10#),
      1481 => to_slv(opcode_type, 16#CD#),
      1482 => to_slv(opcode_type, 16#01#),
      1483 => to_slv(opcode_type, 16#11#),
      1484 => to_slv(opcode_type, 16#07#),
      1485 => to_slv(opcode_type, 16#06#),
      1486 => to_slv(opcode_type, 16#07#),
      1487 => to_slv(opcode_type, 16#0B#),
      1488 => to_slv(opcode_type, 16#10#),
      1489 => to_slv(opcode_type, 16#08#),
      1490 => to_slv(opcode_type, 16#EA#),
      1491 => to_slv(opcode_type, 16#12#),
      1492 => to_slv(opcode_type, 16#06#),
      1493 => to_slv(opcode_type, 16#09#),
      1494 => to_slv(opcode_type, 16#0D#),
      1495 => to_slv(opcode_type, 16#0B#),
      1496 => to_slv(opcode_type, 16#08#),
      1497 => to_slv(opcode_type, 16#0D#),
      1498 => to_slv(opcode_type, 16#0C#),
      1499 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#07#),
      1505 => to_slv(opcode_type, 16#06#),
      1506 => to_slv(opcode_type, 16#02#),
      1507 => to_slv(opcode_type, 16#09#),
      1508 => to_slv(opcode_type, 16#10#),
      1509 => to_slv(opcode_type, 16#10#),
      1510 => to_slv(opcode_type, 16#06#),
      1511 => to_slv(opcode_type, 16#08#),
      1512 => to_slv(opcode_type, 16#10#),
      1513 => to_slv(opcode_type, 16#0D#),
      1514 => to_slv(opcode_type, 16#06#),
      1515 => to_slv(opcode_type, 16#0F#),
      1516 => to_slv(opcode_type, 16#0B#),
      1517 => to_slv(opcode_type, 16#09#),
      1518 => to_slv(opcode_type, 16#08#),
      1519 => to_slv(opcode_type, 16#07#),
      1520 => to_slv(opcode_type, 16#0F#),
      1521 => to_slv(opcode_type, 16#0C#),
      1522 => to_slv(opcode_type, 16#09#),
      1523 => to_slv(opcode_type, 16#11#),
      1524 => to_slv(opcode_type, 16#0F#),
      1525 => to_slv(opcode_type, 16#07#),
      1526 => to_slv(opcode_type, 16#05#),
      1527 => to_slv(opcode_type, 16#11#),
      1528 => to_slv(opcode_type, 16#06#),
      1529 => to_slv(opcode_type, 16#0B#),
      1530 => to_slv(opcode_type, 16#7A#),
      1531 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#07#),
      1537 => to_slv(opcode_type, 16#06#),
      1538 => to_slv(opcode_type, 16#09#),
      1539 => to_slv(opcode_type, 16#04#),
      1540 => to_slv(opcode_type, 16#BE#),
      1541 => to_slv(opcode_type, 16#05#),
      1542 => to_slv(opcode_type, 16#0F#),
      1543 => to_slv(opcode_type, 16#07#),
      1544 => to_slv(opcode_type, 16#05#),
      1545 => to_slv(opcode_type, 16#0F#),
      1546 => to_slv(opcode_type, 16#07#),
      1547 => to_slv(opcode_type, 16#0B#),
      1548 => to_slv(opcode_type, 16#0D#),
      1549 => to_slv(opcode_type, 16#08#),
      1550 => to_slv(opcode_type, 16#09#),
      1551 => to_slv(opcode_type, 16#09#),
      1552 => to_slv(opcode_type, 16#10#),
      1553 => to_slv(opcode_type, 16#0D#),
      1554 => to_slv(opcode_type, 16#04#),
      1555 => to_slv(opcode_type, 16#0A#),
      1556 => to_slv(opcode_type, 16#07#),
      1557 => to_slv(opcode_type, 16#09#),
      1558 => to_slv(opcode_type, 16#0A#),
      1559 => to_slv(opcode_type, 16#10#),
      1560 => to_slv(opcode_type, 16#08#),
      1561 => to_slv(opcode_type, 16#0A#),
      1562 => to_slv(opcode_type, 16#0F#),
      1563 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#09#),
      1569 => to_slv(opcode_type, 16#07#),
      1570 => to_slv(opcode_type, 16#01#),
      1571 => to_slv(opcode_type, 16#09#),
      1572 => to_slv(opcode_type, 16#10#),
      1573 => to_slv(opcode_type, 16#0F#),
      1574 => to_slv(opcode_type, 16#09#),
      1575 => to_slv(opcode_type, 16#03#),
      1576 => to_slv(opcode_type, 16#0D#),
      1577 => to_slv(opcode_type, 16#08#),
      1578 => to_slv(opcode_type, 16#10#),
      1579 => to_slv(opcode_type, 16#10#),
      1580 => to_slv(opcode_type, 16#07#),
      1581 => to_slv(opcode_type, 16#08#),
      1582 => to_slv(opcode_type, 16#07#),
      1583 => to_slv(opcode_type, 16#0A#),
      1584 => to_slv(opcode_type, 16#0C#),
      1585 => to_slv(opcode_type, 16#07#),
      1586 => to_slv(opcode_type, 16#8A#),
      1587 => to_slv(opcode_type, 16#0C#),
      1588 => to_slv(opcode_type, 16#06#),
      1589 => to_slv(opcode_type, 16#09#),
      1590 => to_slv(opcode_type, 16#0A#),
      1591 => to_slv(opcode_type, 16#11#),
      1592 => to_slv(opcode_type, 16#06#),
      1593 => to_slv(opcode_type, 16#0E#),
      1594 => to_slv(opcode_type, 16#0A#),
      1595 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#06#),
      1602 => to_slv(opcode_type, 16#07#),
      1603 => to_slv(opcode_type, 16#02#),
      1604 => to_slv(opcode_type, 16#80#),
      1605 => to_slv(opcode_type, 16#03#),
      1606 => to_slv(opcode_type, 16#0A#),
      1607 => to_slv(opcode_type, 16#06#),
      1608 => to_slv(opcode_type, 16#06#),
      1609 => to_slv(opcode_type, 16#0A#),
      1610 => to_slv(opcode_type, 16#0D#),
      1611 => to_slv(opcode_type, 16#08#),
      1612 => to_slv(opcode_type, 16#0E#),
      1613 => to_slv(opcode_type, 16#0F#),
      1614 => to_slv(opcode_type, 16#06#),
      1615 => to_slv(opcode_type, 16#07#),
      1616 => to_slv(opcode_type, 16#07#),
      1617 => to_slv(opcode_type, 16#0F#),
      1618 => to_slv(opcode_type, 16#0A#),
      1619 => to_slv(opcode_type, 16#04#),
      1620 => to_slv(opcode_type, 16#0D#),
      1621 => to_slv(opcode_type, 16#06#),
      1622 => to_slv(opcode_type, 16#02#),
      1623 => to_slv(opcode_type, 16#10#),
      1624 => to_slv(opcode_type, 16#06#),
      1625 => to_slv(opcode_type, 16#10#),
      1626 => to_slv(opcode_type, 16#0D#),
      1627 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#09#),
      1633 => to_slv(opcode_type, 16#09#),
      1634 => to_slv(opcode_type, 16#01#),
      1635 => to_slv(opcode_type, 16#09#),
      1636 => to_slv(opcode_type, 16#11#),
      1637 => to_slv(opcode_type, 16#0A#),
      1638 => to_slv(opcode_type, 16#08#),
      1639 => to_slv(opcode_type, 16#05#),
      1640 => to_slv(opcode_type, 16#10#),
      1641 => to_slv(opcode_type, 16#07#),
      1642 => to_slv(opcode_type, 16#0A#),
      1643 => to_slv(opcode_type, 16#0B#),
      1644 => to_slv(opcode_type, 16#07#),
      1645 => to_slv(opcode_type, 16#07#),
      1646 => to_slv(opcode_type, 16#06#),
      1647 => to_slv(opcode_type, 16#E9#),
      1648 => to_slv(opcode_type, 16#0B#),
      1649 => to_slv(opcode_type, 16#09#),
      1650 => to_slv(opcode_type, 16#10#),
      1651 => to_slv(opcode_type, 16#1C#),
      1652 => to_slv(opcode_type, 16#07#),
      1653 => to_slv(opcode_type, 16#09#),
      1654 => to_slv(opcode_type, 16#10#),
      1655 => to_slv(opcode_type, 16#10#),
      1656 => to_slv(opcode_type, 16#06#),
      1657 => to_slv(opcode_type, 16#0F#),
      1658 => to_slv(opcode_type, 16#D7#),
      1659 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#07#),
      1665 => to_slv(opcode_type, 16#06#),
      1666 => to_slv(opcode_type, 16#03#),
      1667 => to_slv(opcode_type, 16#05#),
      1668 => to_slv(opcode_type, 16#20#),
      1669 => to_slv(opcode_type, 16#06#),
      1670 => to_slv(opcode_type, 16#06#),
      1671 => to_slv(opcode_type, 16#0E#),
      1672 => to_slv(opcode_type, 16#0A#),
      1673 => to_slv(opcode_type, 16#09#),
      1674 => to_slv(opcode_type, 16#0D#),
      1675 => to_slv(opcode_type, 16#10#),
      1676 => to_slv(opcode_type, 16#09#),
      1677 => to_slv(opcode_type, 16#08#),
      1678 => to_slv(opcode_type, 16#09#),
      1679 => to_slv(opcode_type, 16#0F#),
      1680 => to_slv(opcode_type, 16#0B#),
      1681 => to_slv(opcode_type, 16#07#),
      1682 => to_slv(opcode_type, 16#0F#),
      1683 => to_slv(opcode_type, 16#0D#),
      1684 => to_slv(opcode_type, 16#09#),
      1685 => to_slv(opcode_type, 16#09#),
      1686 => to_slv(opcode_type, 16#0A#),
      1687 => to_slv(opcode_type, 16#0D#),
      1688 => to_slv(opcode_type, 16#08#),
      1689 => to_slv(opcode_type, 16#0D#),
      1690 => to_slv(opcode_type, 16#0B#),
      1691 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#09#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#01#),
      1699 => to_slv(opcode_type, 16#01#),
      1700 => to_slv(opcode_type, 16#0D#),
      1701 => to_slv(opcode_type, 16#08#),
      1702 => to_slv(opcode_type, 16#09#),
      1703 => to_slv(opcode_type, 16#0B#),
      1704 => to_slv(opcode_type, 16#11#),
      1705 => to_slv(opcode_type, 16#07#),
      1706 => to_slv(opcode_type, 16#0C#),
      1707 => to_slv(opcode_type, 16#0D#),
      1708 => to_slv(opcode_type, 16#09#),
      1709 => to_slv(opcode_type, 16#08#),
      1710 => to_slv(opcode_type, 16#09#),
      1711 => to_slv(opcode_type, 16#0E#),
      1712 => to_slv(opcode_type, 16#0E#),
      1713 => to_slv(opcode_type, 16#07#),
      1714 => to_slv(opcode_type, 16#11#),
      1715 => to_slv(opcode_type, 16#0D#),
      1716 => to_slv(opcode_type, 16#08#),
      1717 => to_slv(opcode_type, 16#08#),
      1718 => to_slv(opcode_type, 16#0D#),
      1719 => to_slv(opcode_type, 16#82#),
      1720 => to_slv(opcode_type, 16#09#),
      1721 => to_slv(opcode_type, 16#0D#),
      1722 => to_slv(opcode_type, 16#0C#),
      1723 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#08#),
      1729 => to_slv(opcode_type, 16#08#),
      1730 => to_slv(opcode_type, 16#08#),
      1731 => to_slv(opcode_type, 16#08#),
      1732 => to_slv(opcode_type, 16#10#),
      1733 => to_slv(opcode_type, 16#0F#),
      1734 => to_slv(opcode_type, 16#02#),
      1735 => to_slv(opcode_type, 16#0F#),
      1736 => to_slv(opcode_type, 16#01#),
      1737 => to_slv(opcode_type, 16#06#),
      1738 => to_slv(opcode_type, 16#0C#),
      1739 => to_slv(opcode_type, 16#0D#),
      1740 => to_slv(opcode_type, 16#07#),
      1741 => to_slv(opcode_type, 16#06#),
      1742 => to_slv(opcode_type, 16#08#),
      1743 => to_slv(opcode_type, 16#11#),
      1744 => to_slv(opcode_type, 16#0C#),
      1745 => to_slv(opcode_type, 16#07#),
      1746 => to_slv(opcode_type, 16#0D#),
      1747 => to_slv(opcode_type, 16#0D#),
      1748 => to_slv(opcode_type, 16#08#),
      1749 => to_slv(opcode_type, 16#09#),
      1750 => to_slv(opcode_type, 16#10#),
      1751 => to_slv(opcode_type, 16#0B#),
      1752 => to_slv(opcode_type, 16#09#),
      1753 => to_slv(opcode_type, 16#2C#),
      1754 => to_slv(opcode_type, 16#0C#),
      1755 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#06#),
      1761 => to_slv(opcode_type, 16#06#),
      1762 => to_slv(opcode_type, 16#08#),
      1763 => to_slv(opcode_type, 16#01#),
      1764 => to_slv(opcode_type, 16#0A#),
      1765 => to_slv(opcode_type, 16#06#),
      1766 => to_slv(opcode_type, 16#0D#),
      1767 => to_slv(opcode_type, 16#0E#),
      1768 => to_slv(opcode_type, 16#01#),
      1769 => to_slv(opcode_type, 16#06#),
      1770 => to_slv(opcode_type, 16#10#),
      1771 => to_slv(opcode_type, 16#11#),
      1772 => to_slv(opcode_type, 16#08#),
      1773 => to_slv(opcode_type, 16#08#),
      1774 => to_slv(opcode_type, 16#09#),
      1775 => to_slv(opcode_type, 16#D8#),
      1776 => to_slv(opcode_type, 16#0D#),
      1777 => to_slv(opcode_type, 16#08#),
      1778 => to_slv(opcode_type, 16#0D#),
      1779 => to_slv(opcode_type, 16#0E#),
      1780 => to_slv(opcode_type, 16#09#),
      1781 => to_slv(opcode_type, 16#08#),
      1782 => to_slv(opcode_type, 16#0E#),
      1783 => to_slv(opcode_type, 16#D1#),
      1784 => to_slv(opcode_type, 16#07#),
      1785 => to_slv(opcode_type, 16#0F#),
      1786 => to_slv(opcode_type, 16#0F#),
      1787 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#08#),
      1793 => to_slv(opcode_type, 16#07#),
      1794 => to_slv(opcode_type, 16#01#),
      1795 => to_slv(opcode_type, 16#02#),
      1796 => to_slv(opcode_type, 16#0F#),
      1797 => to_slv(opcode_type, 16#08#),
      1798 => to_slv(opcode_type, 16#09#),
      1799 => to_slv(opcode_type, 16#0F#),
      1800 => to_slv(opcode_type, 16#0D#),
      1801 => to_slv(opcode_type, 16#08#),
      1802 => to_slv(opcode_type, 16#0E#),
      1803 => to_slv(opcode_type, 16#0B#),
      1804 => to_slv(opcode_type, 16#08#),
      1805 => to_slv(opcode_type, 16#07#),
      1806 => to_slv(opcode_type, 16#07#),
      1807 => to_slv(opcode_type, 16#85#),
      1808 => to_slv(opcode_type, 16#0B#),
      1809 => to_slv(opcode_type, 16#07#),
      1810 => to_slv(opcode_type, 16#11#),
      1811 => to_slv(opcode_type, 16#11#),
      1812 => to_slv(opcode_type, 16#08#),
      1813 => to_slv(opcode_type, 16#06#),
      1814 => to_slv(opcode_type, 16#10#),
      1815 => to_slv(opcode_type, 16#0C#),
      1816 => to_slv(opcode_type, 16#07#),
      1817 => to_slv(opcode_type, 16#0A#),
      1818 => to_slv(opcode_type, 16#0A#),
      1819 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#08#),
      1825 => to_slv(opcode_type, 16#08#),
      1826 => to_slv(opcode_type, 16#06#),
      1827 => to_slv(opcode_type, 16#05#),
      1828 => to_slv(opcode_type, 16#0E#),
      1829 => to_slv(opcode_type, 16#05#),
      1830 => to_slv(opcode_type, 16#0B#),
      1831 => to_slv(opcode_type, 16#06#),
      1832 => to_slv(opcode_type, 16#07#),
      1833 => to_slv(opcode_type, 16#0D#),
      1834 => to_slv(opcode_type, 16#0E#),
      1835 => to_slv(opcode_type, 16#02#),
      1836 => to_slv(opcode_type, 16#0F#),
      1837 => to_slv(opcode_type, 16#07#),
      1838 => to_slv(opcode_type, 16#06#),
      1839 => to_slv(opcode_type, 16#04#),
      1840 => to_slv(opcode_type, 16#0E#),
      1841 => to_slv(opcode_type, 16#09#),
      1842 => to_slv(opcode_type, 16#0D#),
      1843 => to_slv(opcode_type, 16#0D#),
      1844 => to_slv(opcode_type, 16#06#),
      1845 => to_slv(opcode_type, 16#08#),
      1846 => to_slv(opcode_type, 16#0F#),
      1847 => to_slv(opcode_type, 16#4A#),
      1848 => to_slv(opcode_type, 16#07#),
      1849 => to_slv(opcode_type, 16#0B#),
      1850 => to_slv(opcode_type, 16#0E#),
      1851 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#08#),
      1857 => to_slv(opcode_type, 16#06#),
      1858 => to_slv(opcode_type, 16#01#),
      1859 => to_slv(opcode_type, 16#07#),
      1860 => to_slv(opcode_type, 16#0C#),
      1861 => to_slv(opcode_type, 16#0F#),
      1862 => to_slv(opcode_type, 16#09#),
      1863 => to_slv(opcode_type, 16#02#),
      1864 => to_slv(opcode_type, 16#0C#),
      1865 => to_slv(opcode_type, 16#07#),
      1866 => to_slv(opcode_type, 16#10#),
      1867 => to_slv(opcode_type, 16#0A#),
      1868 => to_slv(opcode_type, 16#07#),
      1869 => to_slv(opcode_type, 16#08#),
      1870 => to_slv(opcode_type, 16#08#),
      1871 => to_slv(opcode_type, 16#11#),
      1872 => to_slv(opcode_type, 16#0C#),
      1873 => to_slv(opcode_type, 16#06#),
      1874 => to_slv(opcode_type, 16#0B#),
      1875 => to_slv(opcode_type, 16#0A#),
      1876 => to_slv(opcode_type, 16#08#),
      1877 => to_slv(opcode_type, 16#06#),
      1878 => to_slv(opcode_type, 16#0D#),
      1879 => to_slv(opcode_type, 16#0F#),
      1880 => to_slv(opcode_type, 16#07#),
      1881 => to_slv(opcode_type, 16#0F#),
      1882 => to_slv(opcode_type, 16#0C#),
      1883 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#09#),
      1890 => to_slv(opcode_type, 16#09#),
      1891 => to_slv(opcode_type, 16#02#),
      1892 => to_slv(opcode_type, 16#11#),
      1893 => to_slv(opcode_type, 16#08#),
      1894 => to_slv(opcode_type, 16#0A#),
      1895 => to_slv(opcode_type, 16#0B#),
      1896 => to_slv(opcode_type, 16#07#),
      1897 => to_slv(opcode_type, 16#05#),
      1898 => to_slv(opcode_type, 16#0C#),
      1899 => to_slv(opcode_type, 16#09#),
      1900 => to_slv(opcode_type, 16#0C#),
      1901 => to_slv(opcode_type, 16#13#),
      1902 => to_slv(opcode_type, 16#07#),
      1903 => to_slv(opcode_type, 16#09#),
      1904 => to_slv(opcode_type, 16#05#),
      1905 => to_slv(opcode_type, 16#0A#),
      1906 => to_slv(opcode_type, 16#09#),
      1907 => to_slv(opcode_type, 16#0D#),
      1908 => to_slv(opcode_type, 16#0D#),
      1909 => to_slv(opcode_type, 16#06#),
      1910 => to_slv(opcode_type, 16#07#),
      1911 => to_slv(opcode_type, 16#0C#),
      1912 => to_slv(opcode_type, 16#0D#),
      1913 => to_slv(opcode_type, 16#05#),
      1914 => to_slv(opcode_type, 16#10#),
      1915 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#06#),
      1921 => to_slv(opcode_type, 16#08#),
      1922 => to_slv(opcode_type, 16#03#),
      1923 => to_slv(opcode_type, 16#07#),
      1924 => to_slv(opcode_type, 16#87#),
      1925 => to_slv(opcode_type, 16#0C#),
      1926 => to_slv(opcode_type, 16#08#),
      1927 => to_slv(opcode_type, 16#02#),
      1928 => to_slv(opcode_type, 16#F7#),
      1929 => to_slv(opcode_type, 16#07#),
      1930 => to_slv(opcode_type, 16#10#),
      1931 => to_slv(opcode_type, 16#0A#),
      1932 => to_slv(opcode_type, 16#08#),
      1933 => to_slv(opcode_type, 16#06#),
      1934 => to_slv(opcode_type, 16#08#),
      1935 => to_slv(opcode_type, 16#0F#),
      1936 => to_slv(opcode_type, 16#11#),
      1937 => to_slv(opcode_type, 16#07#),
      1938 => to_slv(opcode_type, 16#10#),
      1939 => to_slv(opcode_type, 16#0A#),
      1940 => to_slv(opcode_type, 16#06#),
      1941 => to_slv(opcode_type, 16#09#),
      1942 => to_slv(opcode_type, 16#10#),
      1943 => to_slv(opcode_type, 16#0A#),
      1944 => to_slv(opcode_type, 16#06#),
      1945 => to_slv(opcode_type, 16#0E#),
      1946 => to_slv(opcode_type, 16#44#),
      1947 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#08#),
      1953 => to_slv(opcode_type, 16#08#),
      1954 => to_slv(opcode_type, 16#03#),
      1955 => to_slv(opcode_type, 16#09#),
      1956 => to_slv(opcode_type, 16#0B#),
      1957 => to_slv(opcode_type, 16#11#),
      1958 => to_slv(opcode_type, 16#07#),
      1959 => to_slv(opcode_type, 16#08#),
      1960 => to_slv(opcode_type, 16#10#),
      1961 => to_slv(opcode_type, 16#10#),
      1962 => to_slv(opcode_type, 16#01#),
      1963 => to_slv(opcode_type, 16#0D#),
      1964 => to_slv(opcode_type, 16#06#),
      1965 => to_slv(opcode_type, 16#07#),
      1966 => to_slv(opcode_type, 16#09#),
      1967 => to_slv(opcode_type, 16#0F#),
      1968 => to_slv(opcode_type, 16#0D#),
      1969 => to_slv(opcode_type, 16#08#),
      1970 => to_slv(opcode_type, 16#0F#),
      1971 => to_slv(opcode_type, 16#0B#),
      1972 => to_slv(opcode_type, 16#08#),
      1973 => to_slv(opcode_type, 16#08#),
      1974 => to_slv(opcode_type, 16#0F#),
      1975 => to_slv(opcode_type, 16#11#),
      1976 => to_slv(opcode_type, 16#07#),
      1977 => to_slv(opcode_type, 16#0B#),
      1978 => to_slv(opcode_type, 16#10#),
      1979 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#08#),
      1985 => to_slv(opcode_type, 16#07#),
      1986 => to_slv(opcode_type, 16#07#),
      1987 => to_slv(opcode_type, 16#05#),
      1988 => to_slv(opcode_type, 16#0D#),
      1989 => to_slv(opcode_type, 16#09#),
      1990 => to_slv(opcode_type, 16#7A#),
      1991 => to_slv(opcode_type, 16#0B#),
      1992 => to_slv(opcode_type, 16#05#),
      1993 => to_slv(opcode_type, 16#09#),
      1994 => to_slv(opcode_type, 16#0A#),
      1995 => to_slv(opcode_type, 16#0E#),
      1996 => to_slv(opcode_type, 16#09#),
      1997 => to_slv(opcode_type, 16#06#),
      1998 => to_slv(opcode_type, 16#06#),
      1999 => to_slv(opcode_type, 16#11#),
      2000 => to_slv(opcode_type, 16#0A#),
      2001 => to_slv(opcode_type, 16#09#),
      2002 => to_slv(opcode_type, 16#0F#),
      2003 => to_slv(opcode_type, 16#11#),
      2004 => to_slv(opcode_type, 16#06#),
      2005 => to_slv(opcode_type, 16#09#),
      2006 => to_slv(opcode_type, 16#0B#),
      2007 => to_slv(opcode_type, 16#10#),
      2008 => to_slv(opcode_type, 16#06#),
      2009 => to_slv(opcode_type, 16#0A#),
      2010 => to_slv(opcode_type, 16#11#),
      2011 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#06#),
      2017 => to_slv(opcode_type, 16#09#),
      2018 => to_slv(opcode_type, 16#04#),
      2019 => to_slv(opcode_type, 16#08#),
      2020 => to_slv(opcode_type, 16#0C#),
      2021 => to_slv(opcode_type, 16#0B#),
      2022 => to_slv(opcode_type, 16#06#),
      2023 => to_slv(opcode_type, 16#09#),
      2024 => to_slv(opcode_type, 16#0E#),
      2025 => to_slv(opcode_type, 16#0A#),
      2026 => to_slv(opcode_type, 16#03#),
      2027 => to_slv(opcode_type, 16#0F#),
      2028 => to_slv(opcode_type, 16#06#),
      2029 => to_slv(opcode_type, 16#08#),
      2030 => to_slv(opcode_type, 16#06#),
      2031 => to_slv(opcode_type, 16#31#),
      2032 => to_slv(opcode_type, 16#0B#),
      2033 => to_slv(opcode_type, 16#08#),
      2034 => to_slv(opcode_type, 16#10#),
      2035 => to_slv(opcode_type, 16#11#),
      2036 => to_slv(opcode_type, 16#07#),
      2037 => to_slv(opcode_type, 16#08#),
      2038 => to_slv(opcode_type, 16#0C#),
      2039 => to_slv(opcode_type, 16#0D#),
      2040 => to_slv(opcode_type, 16#07#),
      2041 => to_slv(opcode_type, 16#10#),
      2042 => to_slv(opcode_type, 16#11#),
      2043 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#06#),
      2049 => to_slv(opcode_type, 16#08#),
      2050 => to_slv(opcode_type, 16#05#),
      2051 => to_slv(opcode_type, 16#07#),
      2052 => to_slv(opcode_type, 16#0C#),
      2053 => to_slv(opcode_type, 16#0B#),
      2054 => to_slv(opcode_type, 16#06#),
      2055 => to_slv(opcode_type, 16#04#),
      2056 => to_slv(opcode_type, 16#0C#),
      2057 => to_slv(opcode_type, 16#09#),
      2058 => to_slv(opcode_type, 16#2C#),
      2059 => to_slv(opcode_type, 16#10#),
      2060 => to_slv(opcode_type, 16#06#),
      2061 => to_slv(opcode_type, 16#08#),
      2062 => to_slv(opcode_type, 16#06#),
      2063 => to_slv(opcode_type, 16#0A#),
      2064 => to_slv(opcode_type, 16#0D#),
      2065 => to_slv(opcode_type, 16#08#),
      2066 => to_slv(opcode_type, 16#8E#),
      2067 => to_slv(opcode_type, 16#0F#),
      2068 => to_slv(opcode_type, 16#08#),
      2069 => to_slv(opcode_type, 16#07#),
      2070 => to_slv(opcode_type, 16#0D#),
      2071 => to_slv(opcode_type, 16#0F#),
      2072 => to_slv(opcode_type, 16#07#),
      2073 => to_slv(opcode_type, 16#10#),
      2074 => to_slv(opcode_type, 16#10#),
      2075 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#09#),
      2081 => to_slv(opcode_type, 16#07#),
      2082 => to_slv(opcode_type, 16#08#),
      2083 => to_slv(opcode_type, 16#06#),
      2084 => to_slv(opcode_type, 16#0A#),
      2085 => to_slv(opcode_type, 16#9B#),
      2086 => to_slv(opcode_type, 16#06#),
      2087 => to_slv(opcode_type, 16#11#),
      2088 => to_slv(opcode_type, 16#0B#),
      2089 => to_slv(opcode_type, 16#05#),
      2090 => to_slv(opcode_type, 16#05#),
      2091 => to_slv(opcode_type, 16#11#),
      2092 => to_slv(opcode_type, 16#06#),
      2093 => to_slv(opcode_type, 16#06#),
      2094 => to_slv(opcode_type, 16#08#),
      2095 => to_slv(opcode_type, 16#0C#),
      2096 => to_slv(opcode_type, 16#0C#),
      2097 => to_slv(opcode_type, 16#08#),
      2098 => to_slv(opcode_type, 16#5E#),
      2099 => to_slv(opcode_type, 16#0B#),
      2100 => to_slv(opcode_type, 16#09#),
      2101 => to_slv(opcode_type, 16#06#),
      2102 => to_slv(opcode_type, 16#11#),
      2103 => to_slv(opcode_type, 16#0D#),
      2104 => to_slv(opcode_type, 16#09#),
      2105 => to_slv(opcode_type, 16#0D#),
      2106 => to_slv(opcode_type, 16#0E#),
      2107 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#09#),
      2113 => to_slv(opcode_type, 16#09#),
      2114 => to_slv(opcode_type, 16#06#),
      2115 => to_slv(opcode_type, 16#09#),
      2116 => to_slv(opcode_type, 16#0A#),
      2117 => to_slv(opcode_type, 16#10#),
      2118 => to_slv(opcode_type, 16#05#),
      2119 => to_slv(opcode_type, 16#0E#),
      2120 => to_slv(opcode_type, 16#07#),
      2121 => to_slv(opcode_type, 16#01#),
      2122 => to_slv(opcode_type, 16#0A#),
      2123 => to_slv(opcode_type, 16#04#),
      2124 => to_slv(opcode_type, 16#0E#),
      2125 => to_slv(opcode_type, 16#08#),
      2126 => to_slv(opcode_type, 16#09#),
      2127 => to_slv(opcode_type, 16#08#),
      2128 => to_slv(opcode_type, 16#0F#),
      2129 => to_slv(opcode_type, 16#0E#),
      2130 => to_slv(opcode_type, 16#09#),
      2131 => to_slv(opcode_type, 16#0C#),
      2132 => to_slv(opcode_type, 16#0D#),
      2133 => to_slv(opcode_type, 16#07#),
      2134 => to_slv(opcode_type, 16#06#),
      2135 => to_slv(opcode_type, 16#0C#),
      2136 => to_slv(opcode_type, 16#0C#),
      2137 => to_slv(opcode_type, 16#04#),
      2138 => to_slv(opcode_type, 16#10#),
      2139 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#07#),
      2145 => to_slv(opcode_type, 16#07#),
      2146 => to_slv(opcode_type, 16#01#),
      2147 => to_slv(opcode_type, 16#09#),
      2148 => to_slv(opcode_type, 16#0E#),
      2149 => to_slv(opcode_type, 16#0F#),
      2150 => to_slv(opcode_type, 16#07#),
      2151 => to_slv(opcode_type, 16#08#),
      2152 => to_slv(opcode_type, 16#0E#),
      2153 => to_slv(opcode_type, 16#0E#),
      2154 => to_slv(opcode_type, 16#06#),
      2155 => to_slv(opcode_type, 16#0A#),
      2156 => to_slv(opcode_type, 16#0F#),
      2157 => to_slv(opcode_type, 16#06#),
      2158 => to_slv(opcode_type, 16#08#),
      2159 => to_slv(opcode_type, 16#01#),
      2160 => to_slv(opcode_type, 16#0D#),
      2161 => to_slv(opcode_type, 16#09#),
      2162 => to_slv(opcode_type, 16#0A#),
      2163 => to_slv(opcode_type, 16#0F#),
      2164 => to_slv(opcode_type, 16#06#),
      2165 => to_slv(opcode_type, 16#09#),
      2166 => to_slv(opcode_type, 16#0A#),
      2167 => to_slv(opcode_type, 16#0A#),
      2168 => to_slv(opcode_type, 16#06#),
      2169 => to_slv(opcode_type, 16#0B#),
      2170 => to_slv(opcode_type, 16#0C#),
      2171 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#09#),
      2177 => to_slv(opcode_type, 16#07#),
      2178 => to_slv(opcode_type, 16#06#),
      2179 => to_slv(opcode_type, 16#08#),
      2180 => to_slv(opcode_type, 16#0C#),
      2181 => to_slv(opcode_type, 16#0E#),
      2182 => to_slv(opcode_type, 16#01#),
      2183 => to_slv(opcode_type, 16#11#),
      2184 => to_slv(opcode_type, 16#08#),
      2185 => to_slv(opcode_type, 16#08#),
      2186 => to_slv(opcode_type, 16#F4#),
      2187 => to_slv(opcode_type, 16#10#),
      2188 => to_slv(opcode_type, 16#04#),
      2189 => to_slv(opcode_type, 16#0A#),
      2190 => to_slv(opcode_type, 16#07#),
      2191 => to_slv(opcode_type, 16#06#),
      2192 => to_slv(opcode_type, 16#01#),
      2193 => to_slv(opcode_type, 16#11#),
      2194 => to_slv(opcode_type, 16#03#),
      2195 => to_slv(opcode_type, 16#23#),
      2196 => to_slv(opcode_type, 16#07#),
      2197 => to_slv(opcode_type, 16#08#),
      2198 => to_slv(opcode_type, 16#0B#),
      2199 => to_slv(opcode_type, 16#0E#),
      2200 => to_slv(opcode_type, 16#07#),
      2201 => to_slv(opcode_type, 16#0A#),
      2202 => to_slv(opcode_type, 16#0B#),
      2203 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#07#),
      2209 => to_slv(opcode_type, 16#07#),
      2210 => to_slv(opcode_type, 16#07#),
      2211 => to_slv(opcode_type, 16#05#),
      2212 => to_slv(opcode_type, 16#0E#),
      2213 => to_slv(opcode_type, 16#02#),
      2214 => to_slv(opcode_type, 16#0A#),
      2215 => to_slv(opcode_type, 16#09#),
      2216 => to_slv(opcode_type, 16#08#),
      2217 => to_slv(opcode_type, 16#0A#),
      2218 => to_slv(opcode_type, 16#0B#),
      2219 => to_slv(opcode_type, 16#07#),
      2220 => to_slv(opcode_type, 16#10#),
      2221 => to_slv(opcode_type, 16#0B#),
      2222 => to_slv(opcode_type, 16#09#),
      2223 => to_slv(opcode_type, 16#08#),
      2224 => to_slv(opcode_type, 16#09#),
      2225 => to_slv(opcode_type, 16#10#),
      2226 => to_slv(opcode_type, 16#0A#),
      2227 => to_slv(opcode_type, 16#06#),
      2228 => to_slv(opcode_type, 16#BA#),
      2229 => to_slv(opcode_type, 16#10#),
      2230 => to_slv(opcode_type, 16#09#),
      2231 => to_slv(opcode_type, 16#05#),
      2232 => to_slv(opcode_type, 16#CB#),
      2233 => to_slv(opcode_type, 16#05#),
      2234 => to_slv(opcode_type, 16#0C#),
      2235 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#08#),
      2242 => to_slv(opcode_type, 16#04#),
      2243 => to_slv(opcode_type, 16#06#),
      2244 => to_slv(opcode_type, 16#0C#),
      2245 => to_slv(opcode_type, 16#0B#),
      2246 => to_slv(opcode_type, 16#07#),
      2247 => to_slv(opcode_type, 16#03#),
      2248 => to_slv(opcode_type, 16#11#),
      2249 => to_slv(opcode_type, 16#09#),
      2250 => to_slv(opcode_type, 16#0A#),
      2251 => to_slv(opcode_type, 16#0D#),
      2252 => to_slv(opcode_type, 16#07#),
      2253 => to_slv(opcode_type, 16#08#),
      2254 => to_slv(opcode_type, 16#08#),
      2255 => to_slv(opcode_type, 16#0C#),
      2256 => to_slv(opcode_type, 16#0D#),
      2257 => to_slv(opcode_type, 16#07#),
      2258 => to_slv(opcode_type, 16#0E#),
      2259 => to_slv(opcode_type, 16#0A#),
      2260 => to_slv(opcode_type, 16#07#),
      2261 => to_slv(opcode_type, 16#07#),
      2262 => to_slv(opcode_type, 16#11#),
      2263 => to_slv(opcode_type, 16#DF#),
      2264 => to_slv(opcode_type, 16#06#),
      2265 => to_slv(opcode_type, 16#0B#),
      2266 => to_slv(opcode_type, 16#0D#),
      2267 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#06#),
      2273 => to_slv(opcode_type, 16#07#),
      2274 => to_slv(opcode_type, 16#06#),
      2275 => to_slv(opcode_type, 16#05#),
      2276 => to_slv(opcode_type, 16#D3#),
      2277 => to_slv(opcode_type, 16#07#),
      2278 => to_slv(opcode_type, 16#0F#),
      2279 => to_slv(opcode_type, 16#11#),
      2280 => to_slv(opcode_type, 16#02#),
      2281 => to_slv(opcode_type, 16#06#),
      2282 => to_slv(opcode_type, 16#0A#),
      2283 => to_slv(opcode_type, 16#0A#),
      2284 => to_slv(opcode_type, 16#06#),
      2285 => to_slv(opcode_type, 16#07#),
      2286 => to_slv(opcode_type, 16#07#),
      2287 => to_slv(opcode_type, 16#0A#),
      2288 => to_slv(opcode_type, 16#1F#),
      2289 => to_slv(opcode_type, 16#09#),
      2290 => to_slv(opcode_type, 16#10#),
      2291 => to_slv(opcode_type, 16#11#),
      2292 => to_slv(opcode_type, 16#07#),
      2293 => to_slv(opcode_type, 16#07#),
      2294 => to_slv(opcode_type, 16#7B#),
      2295 => to_slv(opcode_type, 16#10#),
      2296 => to_slv(opcode_type, 16#09#),
      2297 => to_slv(opcode_type, 16#0A#),
      2298 => to_slv(opcode_type, 16#0B#),
      2299 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#07#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#07#),
      2307 => to_slv(opcode_type, 16#08#),
      2308 => to_slv(opcode_type, 16#0B#),
      2309 => to_slv(opcode_type, 16#10#),
      2310 => to_slv(opcode_type, 16#01#),
      2311 => to_slv(opcode_type, 16#11#),
      2312 => to_slv(opcode_type, 16#04#),
      2313 => to_slv(opcode_type, 16#07#),
      2314 => to_slv(opcode_type, 16#0B#),
      2315 => to_slv(opcode_type, 16#0B#),
      2316 => to_slv(opcode_type, 16#06#),
      2317 => to_slv(opcode_type, 16#08#),
      2318 => to_slv(opcode_type, 16#07#),
      2319 => to_slv(opcode_type, 16#57#),
      2320 => to_slv(opcode_type, 16#0F#),
      2321 => to_slv(opcode_type, 16#09#),
      2322 => to_slv(opcode_type, 16#0E#),
      2323 => to_slv(opcode_type, 16#0D#),
      2324 => to_slv(opcode_type, 16#07#),
      2325 => to_slv(opcode_type, 16#08#),
      2326 => to_slv(opcode_type, 16#0B#),
      2327 => to_slv(opcode_type, 16#0B#),
      2328 => to_slv(opcode_type, 16#07#),
      2329 => to_slv(opcode_type, 16#11#),
      2330 => to_slv(opcode_type, 16#E8#),
      2331 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#07#),
      2337 => to_slv(opcode_type, 16#07#),
      2338 => to_slv(opcode_type, 16#06#),
      2339 => to_slv(opcode_type, 16#03#),
      2340 => to_slv(opcode_type, 16#0F#),
      2341 => to_slv(opcode_type, 16#04#),
      2342 => to_slv(opcode_type, 16#0C#),
      2343 => to_slv(opcode_type, 16#07#),
      2344 => to_slv(opcode_type, 16#08#),
      2345 => to_slv(opcode_type, 16#0F#),
      2346 => to_slv(opcode_type, 16#F2#),
      2347 => to_slv(opcode_type, 16#09#),
      2348 => to_slv(opcode_type, 16#0A#),
      2349 => to_slv(opcode_type, 16#CD#),
      2350 => to_slv(opcode_type, 16#07#),
      2351 => to_slv(opcode_type, 16#09#),
      2352 => to_slv(opcode_type, 16#06#),
      2353 => to_slv(opcode_type, 16#0E#),
      2354 => to_slv(opcode_type, 16#11#),
      2355 => to_slv(opcode_type, 16#02#),
      2356 => to_slv(opcode_type, 16#B6#),
      2357 => to_slv(opcode_type, 16#06#),
      2358 => to_slv(opcode_type, 16#01#),
      2359 => to_slv(opcode_type, 16#0C#),
      2360 => to_slv(opcode_type, 16#06#),
      2361 => to_slv(opcode_type, 16#11#),
      2362 => to_slv(opcode_type, 16#EB#),
      2363 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#06#),
      2369 => to_slv(opcode_type, 16#06#),
      2370 => to_slv(opcode_type, 16#05#),
      2371 => to_slv(opcode_type, 16#08#),
      2372 => to_slv(opcode_type, 16#0D#),
      2373 => to_slv(opcode_type, 16#0D#),
      2374 => to_slv(opcode_type, 16#06#),
      2375 => to_slv(opcode_type, 16#04#),
      2376 => to_slv(opcode_type, 16#0B#),
      2377 => to_slv(opcode_type, 16#07#),
      2378 => to_slv(opcode_type, 16#0D#),
      2379 => to_slv(opcode_type, 16#11#),
      2380 => to_slv(opcode_type, 16#08#),
      2381 => to_slv(opcode_type, 16#07#),
      2382 => to_slv(opcode_type, 16#08#),
      2383 => to_slv(opcode_type, 16#0B#),
      2384 => to_slv(opcode_type, 16#11#),
      2385 => to_slv(opcode_type, 16#08#),
      2386 => to_slv(opcode_type, 16#0F#),
      2387 => to_slv(opcode_type, 16#0F#),
      2388 => to_slv(opcode_type, 16#09#),
      2389 => to_slv(opcode_type, 16#06#),
      2390 => to_slv(opcode_type, 16#11#),
      2391 => to_slv(opcode_type, 16#0F#),
      2392 => to_slv(opcode_type, 16#09#),
      2393 => to_slv(opcode_type, 16#C0#),
      2394 => to_slv(opcode_type, 16#0B#),
      2395 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#06#),
      2402 => to_slv(opcode_type, 16#09#),
      2403 => to_slv(opcode_type, 16#03#),
      2404 => to_slv(opcode_type, 16#0C#),
      2405 => to_slv(opcode_type, 16#09#),
      2406 => to_slv(opcode_type, 16#0F#),
      2407 => to_slv(opcode_type, 16#0C#),
      2408 => to_slv(opcode_type, 16#08#),
      2409 => to_slv(opcode_type, 16#09#),
      2410 => to_slv(opcode_type, 16#0A#),
      2411 => to_slv(opcode_type, 16#0D#),
      2412 => to_slv(opcode_type, 16#01#),
      2413 => to_slv(opcode_type, 16#10#),
      2414 => to_slv(opcode_type, 16#06#),
      2415 => to_slv(opcode_type, 16#09#),
      2416 => to_slv(opcode_type, 16#07#),
      2417 => to_slv(opcode_type, 16#0F#),
      2418 => to_slv(opcode_type, 16#0E#),
      2419 => to_slv(opcode_type, 16#09#),
      2420 => to_slv(opcode_type, 16#0D#),
      2421 => to_slv(opcode_type, 16#C4#),
      2422 => to_slv(opcode_type, 16#08#),
      2423 => to_slv(opcode_type, 16#09#),
      2424 => to_slv(opcode_type, 16#0B#),
      2425 => to_slv(opcode_type, 16#64#),
      2426 => to_slv(opcode_type, 16#0C#),
      2427 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#09#),
      2433 => to_slv(opcode_type, 16#09#),
      2434 => to_slv(opcode_type, 16#05#),
      2435 => to_slv(opcode_type, 16#03#),
      2436 => to_slv(opcode_type, 16#0E#),
      2437 => to_slv(opcode_type, 16#09#),
      2438 => to_slv(opcode_type, 16#09#),
      2439 => to_slv(opcode_type, 16#0D#),
      2440 => to_slv(opcode_type, 16#0F#),
      2441 => to_slv(opcode_type, 16#06#),
      2442 => to_slv(opcode_type, 16#11#),
      2443 => to_slv(opcode_type, 16#C4#),
      2444 => to_slv(opcode_type, 16#09#),
      2445 => to_slv(opcode_type, 16#08#),
      2446 => to_slv(opcode_type, 16#08#),
      2447 => to_slv(opcode_type, 16#0B#),
      2448 => to_slv(opcode_type, 16#0F#),
      2449 => to_slv(opcode_type, 16#09#),
      2450 => to_slv(opcode_type, 16#0B#),
      2451 => to_slv(opcode_type, 16#0C#),
      2452 => to_slv(opcode_type, 16#08#),
      2453 => to_slv(opcode_type, 16#06#),
      2454 => to_slv(opcode_type, 16#10#),
      2455 => to_slv(opcode_type, 16#0B#),
      2456 => to_slv(opcode_type, 16#07#),
      2457 => to_slv(opcode_type, 16#0D#),
      2458 => to_slv(opcode_type, 16#0A#),
      2459 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#06#),
      2465 => to_slv(opcode_type, 16#08#),
      2466 => to_slv(opcode_type, 16#04#),
      2467 => to_slv(opcode_type, 16#09#),
      2468 => to_slv(opcode_type, 16#0C#),
      2469 => to_slv(opcode_type, 16#0D#),
      2470 => to_slv(opcode_type, 16#08#),
      2471 => to_slv(opcode_type, 16#07#),
      2472 => to_slv(opcode_type, 16#0E#),
      2473 => to_slv(opcode_type, 16#0B#),
      2474 => to_slv(opcode_type, 16#02#),
      2475 => to_slv(opcode_type, 16#0C#),
      2476 => to_slv(opcode_type, 16#08#),
      2477 => to_slv(opcode_type, 16#06#),
      2478 => to_slv(opcode_type, 16#07#),
      2479 => to_slv(opcode_type, 16#0F#),
      2480 => to_slv(opcode_type, 16#BF#),
      2481 => to_slv(opcode_type, 16#06#),
      2482 => to_slv(opcode_type, 16#0F#),
      2483 => to_slv(opcode_type, 16#19#),
      2484 => to_slv(opcode_type, 16#08#),
      2485 => to_slv(opcode_type, 16#09#),
      2486 => to_slv(opcode_type, 16#11#),
      2487 => to_slv(opcode_type, 16#11#),
      2488 => to_slv(opcode_type, 16#07#),
      2489 => to_slv(opcode_type, 16#0F#),
      2490 => to_slv(opcode_type, 16#0E#),
      2491 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#08#),
      2497 => to_slv(opcode_type, 16#09#),
      2498 => to_slv(opcode_type, 16#03#),
      2499 => to_slv(opcode_type, 16#09#),
      2500 => to_slv(opcode_type, 16#11#),
      2501 => to_slv(opcode_type, 16#0D#),
      2502 => to_slv(opcode_type, 16#07#),
      2503 => to_slv(opcode_type, 16#05#),
      2504 => to_slv(opcode_type, 16#0C#),
      2505 => to_slv(opcode_type, 16#07#),
      2506 => to_slv(opcode_type, 16#11#),
      2507 => to_slv(opcode_type, 16#58#),
      2508 => to_slv(opcode_type, 16#06#),
      2509 => to_slv(opcode_type, 16#09#),
      2510 => to_slv(opcode_type, 16#09#),
      2511 => to_slv(opcode_type, 16#10#),
      2512 => to_slv(opcode_type, 16#0D#),
      2513 => to_slv(opcode_type, 16#08#),
      2514 => to_slv(opcode_type, 16#0F#),
      2515 => to_slv(opcode_type, 16#10#),
      2516 => to_slv(opcode_type, 16#09#),
      2517 => to_slv(opcode_type, 16#08#),
      2518 => to_slv(opcode_type, 16#0D#),
      2519 => to_slv(opcode_type, 16#0B#),
      2520 => to_slv(opcode_type, 16#07#),
      2521 => to_slv(opcode_type, 16#0F#),
      2522 => to_slv(opcode_type, 16#11#),
      2523 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#06#),
      2529 => to_slv(opcode_type, 16#08#),
      2530 => to_slv(opcode_type, 16#01#),
      2531 => to_slv(opcode_type, 16#02#),
      2532 => to_slv(opcode_type, 16#0C#),
      2533 => to_slv(opcode_type, 16#09#),
      2534 => to_slv(opcode_type, 16#09#),
      2535 => to_slv(opcode_type, 16#0E#),
      2536 => to_slv(opcode_type, 16#10#),
      2537 => to_slv(opcode_type, 16#07#),
      2538 => to_slv(opcode_type, 16#0D#),
      2539 => to_slv(opcode_type, 16#0B#),
      2540 => to_slv(opcode_type, 16#09#),
      2541 => to_slv(opcode_type, 16#09#),
      2542 => to_slv(opcode_type, 16#09#),
      2543 => to_slv(opcode_type, 16#0E#),
      2544 => to_slv(opcode_type, 16#10#),
      2545 => to_slv(opcode_type, 16#09#),
      2546 => to_slv(opcode_type, 16#10#),
      2547 => to_slv(opcode_type, 16#0A#),
      2548 => to_slv(opcode_type, 16#08#),
      2549 => to_slv(opcode_type, 16#07#),
      2550 => to_slv(opcode_type, 16#10#),
      2551 => to_slv(opcode_type, 16#0C#),
      2552 => to_slv(opcode_type, 16#07#),
      2553 => to_slv(opcode_type, 16#0F#),
      2554 => to_slv(opcode_type, 16#0D#),
      2555 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#08#),
      2561 => to_slv(opcode_type, 16#06#),
      2562 => to_slv(opcode_type, 16#05#),
      2563 => to_slv(opcode_type, 16#03#),
      2564 => to_slv(opcode_type, 16#0B#),
      2565 => to_slv(opcode_type, 16#07#),
      2566 => to_slv(opcode_type, 16#08#),
      2567 => to_slv(opcode_type, 16#0B#),
      2568 => to_slv(opcode_type, 16#0C#),
      2569 => to_slv(opcode_type, 16#06#),
      2570 => to_slv(opcode_type, 16#1F#),
      2571 => to_slv(opcode_type, 16#AC#),
      2572 => to_slv(opcode_type, 16#07#),
      2573 => to_slv(opcode_type, 16#06#),
      2574 => to_slv(opcode_type, 16#07#),
      2575 => to_slv(opcode_type, 16#B0#),
      2576 => to_slv(opcode_type, 16#0C#),
      2577 => to_slv(opcode_type, 16#09#),
      2578 => to_slv(opcode_type, 16#42#),
      2579 => to_slv(opcode_type, 16#0F#),
      2580 => to_slv(opcode_type, 16#08#),
      2581 => to_slv(opcode_type, 16#09#),
      2582 => to_slv(opcode_type, 16#0E#),
      2583 => to_slv(opcode_type, 16#0C#),
      2584 => to_slv(opcode_type, 16#09#),
      2585 => to_slv(opcode_type, 16#10#),
      2586 => to_slv(opcode_type, 16#11#),
      2587 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#07#),
      2593 => to_slv(opcode_type, 16#07#),
      2594 => to_slv(opcode_type, 16#05#),
      2595 => to_slv(opcode_type, 16#04#),
      2596 => to_slv(opcode_type, 16#10#),
      2597 => to_slv(opcode_type, 16#09#),
      2598 => to_slv(opcode_type, 16#07#),
      2599 => to_slv(opcode_type, 16#0A#),
      2600 => to_slv(opcode_type, 16#21#),
      2601 => to_slv(opcode_type, 16#07#),
      2602 => to_slv(opcode_type, 16#0F#),
      2603 => to_slv(opcode_type, 16#0F#),
      2604 => to_slv(opcode_type, 16#06#),
      2605 => to_slv(opcode_type, 16#08#),
      2606 => to_slv(opcode_type, 16#07#),
      2607 => to_slv(opcode_type, 16#9A#),
      2608 => to_slv(opcode_type, 16#C5#),
      2609 => to_slv(opcode_type, 16#09#),
      2610 => to_slv(opcode_type, 16#11#),
      2611 => to_slv(opcode_type, 16#0E#),
      2612 => to_slv(opcode_type, 16#07#),
      2613 => to_slv(opcode_type, 16#08#),
      2614 => to_slv(opcode_type, 16#11#),
      2615 => to_slv(opcode_type, 16#10#),
      2616 => to_slv(opcode_type, 16#08#),
      2617 => to_slv(opcode_type, 16#0A#),
      2618 => to_slv(opcode_type, 16#10#),
      2619 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#06#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#09#),
      2627 => to_slv(opcode_type, 16#09#),
      2628 => to_slv(opcode_type, 16#0D#),
      2629 => to_slv(opcode_type, 16#10#),
      2630 => to_slv(opcode_type, 16#05#),
      2631 => to_slv(opcode_type, 16#10#),
      2632 => to_slv(opcode_type, 16#02#),
      2633 => to_slv(opcode_type, 16#07#),
      2634 => to_slv(opcode_type, 16#0C#),
      2635 => to_slv(opcode_type, 16#0F#),
      2636 => to_slv(opcode_type, 16#09#),
      2637 => to_slv(opcode_type, 16#06#),
      2638 => to_slv(opcode_type, 16#07#),
      2639 => to_slv(opcode_type, 16#0C#),
      2640 => to_slv(opcode_type, 16#0A#),
      2641 => to_slv(opcode_type, 16#06#),
      2642 => to_slv(opcode_type, 16#0F#),
      2643 => to_slv(opcode_type, 16#37#),
      2644 => to_slv(opcode_type, 16#09#),
      2645 => to_slv(opcode_type, 16#07#),
      2646 => to_slv(opcode_type, 16#0A#),
      2647 => to_slv(opcode_type, 16#11#),
      2648 => to_slv(opcode_type, 16#07#),
      2649 => to_slv(opcode_type, 16#10#),
      2650 => to_slv(opcode_type, 16#95#),
      2651 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#07#),
      2657 => to_slv(opcode_type, 16#07#),
      2658 => to_slv(opcode_type, 16#09#),
      2659 => to_slv(opcode_type, 16#02#),
      2660 => to_slv(opcode_type, 16#0D#),
      2661 => to_slv(opcode_type, 16#08#),
      2662 => to_slv(opcode_type, 16#0A#),
      2663 => to_slv(opcode_type, 16#0E#),
      2664 => to_slv(opcode_type, 16#04#),
      2665 => to_slv(opcode_type, 16#09#),
      2666 => to_slv(opcode_type, 16#0D#),
      2667 => to_slv(opcode_type, 16#0B#),
      2668 => to_slv(opcode_type, 16#09#),
      2669 => to_slv(opcode_type, 16#07#),
      2670 => to_slv(opcode_type, 16#07#),
      2671 => to_slv(opcode_type, 16#0E#),
      2672 => to_slv(opcode_type, 16#A0#),
      2673 => to_slv(opcode_type, 16#09#),
      2674 => to_slv(opcode_type, 16#0B#),
      2675 => to_slv(opcode_type, 16#0F#),
      2676 => to_slv(opcode_type, 16#08#),
      2677 => to_slv(opcode_type, 16#08#),
      2678 => to_slv(opcode_type, 16#11#),
      2679 => to_slv(opcode_type, 16#11#),
      2680 => to_slv(opcode_type, 16#09#),
      2681 => to_slv(opcode_type, 16#0F#),
      2682 => to_slv(opcode_type, 16#10#),
      2683 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#08#),
      2689 => to_slv(opcode_type, 16#06#),
      2690 => to_slv(opcode_type, 16#02#),
      2691 => to_slv(opcode_type, 16#07#),
      2692 => to_slv(opcode_type, 16#0E#),
      2693 => to_slv(opcode_type, 16#0F#),
      2694 => to_slv(opcode_type, 16#09#),
      2695 => to_slv(opcode_type, 16#07#),
      2696 => to_slv(opcode_type, 16#10#),
      2697 => to_slv(opcode_type, 16#0B#),
      2698 => to_slv(opcode_type, 16#03#),
      2699 => to_slv(opcode_type, 16#0A#),
      2700 => to_slv(opcode_type, 16#08#),
      2701 => to_slv(opcode_type, 16#09#),
      2702 => to_slv(opcode_type, 16#07#),
      2703 => to_slv(opcode_type, 16#0E#),
      2704 => to_slv(opcode_type, 16#10#),
      2705 => to_slv(opcode_type, 16#09#),
      2706 => to_slv(opcode_type, 16#0A#),
      2707 => to_slv(opcode_type, 16#0F#),
      2708 => to_slv(opcode_type, 16#09#),
      2709 => to_slv(opcode_type, 16#09#),
      2710 => to_slv(opcode_type, 16#11#),
      2711 => to_slv(opcode_type, 16#DB#),
      2712 => to_slv(opcode_type, 16#09#),
      2713 => to_slv(opcode_type, 16#0C#),
      2714 => to_slv(opcode_type, 16#0E#),
      2715 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#07#),
      2721 => to_slv(opcode_type, 16#08#),
      2722 => to_slv(opcode_type, 16#01#),
      2723 => to_slv(opcode_type, 16#09#),
      2724 => to_slv(opcode_type, 16#0D#),
      2725 => to_slv(opcode_type, 16#10#),
      2726 => to_slv(opcode_type, 16#08#),
      2727 => to_slv(opcode_type, 16#09#),
      2728 => to_slv(opcode_type, 16#0E#),
      2729 => to_slv(opcode_type, 16#0D#),
      2730 => to_slv(opcode_type, 16#07#),
      2731 => to_slv(opcode_type, 16#11#),
      2732 => to_slv(opcode_type, 16#11#),
      2733 => to_slv(opcode_type, 16#09#),
      2734 => to_slv(opcode_type, 16#07#),
      2735 => to_slv(opcode_type, 16#03#),
      2736 => to_slv(opcode_type, 16#10#),
      2737 => to_slv(opcode_type, 16#08#),
      2738 => to_slv(opcode_type, 16#0B#),
      2739 => to_slv(opcode_type, 16#0B#),
      2740 => to_slv(opcode_type, 16#06#),
      2741 => to_slv(opcode_type, 16#09#),
      2742 => to_slv(opcode_type, 16#0E#),
      2743 => to_slv(opcode_type, 16#0B#),
      2744 => to_slv(opcode_type, 16#09#),
      2745 => to_slv(opcode_type, 16#0C#),
      2746 => to_slv(opcode_type, 16#0F#),
      2747 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#08#),
      2753 => to_slv(opcode_type, 16#09#),
      2754 => to_slv(opcode_type, 16#08#),
      2755 => to_slv(opcode_type, 16#09#),
      2756 => to_slv(opcode_type, 16#0A#),
      2757 => to_slv(opcode_type, 16#11#),
      2758 => to_slv(opcode_type, 16#02#),
      2759 => to_slv(opcode_type, 16#0E#),
      2760 => to_slv(opcode_type, 16#04#),
      2761 => to_slv(opcode_type, 16#08#),
      2762 => to_slv(opcode_type, 16#0F#),
      2763 => to_slv(opcode_type, 16#0D#),
      2764 => to_slv(opcode_type, 16#07#),
      2765 => to_slv(opcode_type, 16#07#),
      2766 => to_slv(opcode_type, 16#09#),
      2767 => to_slv(opcode_type, 16#0D#),
      2768 => to_slv(opcode_type, 16#0A#),
      2769 => to_slv(opcode_type, 16#09#),
      2770 => to_slv(opcode_type, 16#0A#),
      2771 => to_slv(opcode_type, 16#0B#),
      2772 => to_slv(opcode_type, 16#06#),
      2773 => to_slv(opcode_type, 16#07#),
      2774 => to_slv(opcode_type, 16#0C#),
      2775 => to_slv(opcode_type, 16#0B#),
      2776 => to_slv(opcode_type, 16#07#),
      2777 => to_slv(opcode_type, 16#11#),
      2778 => to_slv(opcode_type, 16#0C#),
      2779 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#08#),
      2785 => to_slv(opcode_type, 16#08#),
      2786 => to_slv(opcode_type, 16#05#),
      2787 => to_slv(opcode_type, 16#03#),
      2788 => to_slv(opcode_type, 16#0B#),
      2789 => to_slv(opcode_type, 16#07#),
      2790 => to_slv(opcode_type, 16#09#),
      2791 => to_slv(opcode_type, 16#10#),
      2792 => to_slv(opcode_type, 16#10#),
      2793 => to_slv(opcode_type, 16#07#),
      2794 => to_slv(opcode_type, 16#11#),
      2795 => to_slv(opcode_type, 16#89#),
      2796 => to_slv(opcode_type, 16#06#),
      2797 => to_slv(opcode_type, 16#09#),
      2798 => to_slv(opcode_type, 16#07#),
      2799 => to_slv(opcode_type, 16#10#),
      2800 => to_slv(opcode_type, 16#0A#),
      2801 => to_slv(opcode_type, 16#09#),
      2802 => to_slv(opcode_type, 16#0E#),
      2803 => to_slv(opcode_type, 16#0E#),
      2804 => to_slv(opcode_type, 16#06#),
      2805 => to_slv(opcode_type, 16#07#),
      2806 => to_slv(opcode_type, 16#22#),
      2807 => to_slv(opcode_type, 16#10#),
      2808 => to_slv(opcode_type, 16#06#),
      2809 => to_slv(opcode_type, 16#0B#),
      2810 => to_slv(opcode_type, 16#11#),
      2811 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#09#),
      2817 => to_slv(opcode_type, 16#08#),
      2818 => to_slv(opcode_type, 16#01#),
      2819 => to_slv(opcode_type, 16#07#),
      2820 => to_slv(opcode_type, 16#0B#),
      2821 => to_slv(opcode_type, 16#0E#),
      2822 => to_slv(opcode_type, 16#06#),
      2823 => to_slv(opcode_type, 16#07#),
      2824 => to_slv(opcode_type, 16#0A#),
      2825 => to_slv(opcode_type, 16#0F#),
      2826 => to_slv(opcode_type, 16#06#),
      2827 => to_slv(opcode_type, 16#0D#),
      2828 => to_slv(opcode_type, 16#0A#),
      2829 => to_slv(opcode_type, 16#08#),
      2830 => to_slv(opcode_type, 16#09#),
      2831 => to_slv(opcode_type, 16#02#),
      2832 => to_slv(opcode_type, 16#0D#),
      2833 => to_slv(opcode_type, 16#09#),
      2834 => to_slv(opcode_type, 16#57#),
      2835 => to_slv(opcode_type, 16#0B#),
      2836 => to_slv(opcode_type, 16#07#),
      2837 => to_slv(opcode_type, 16#09#),
      2838 => to_slv(opcode_type, 16#0B#),
      2839 => to_slv(opcode_type, 16#10#),
      2840 => to_slv(opcode_type, 16#08#),
      2841 => to_slv(opcode_type, 16#0B#),
      2842 => to_slv(opcode_type, 16#10#),
      2843 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#06#),
      2849 => to_slv(opcode_type, 16#06#),
      2850 => to_slv(opcode_type, 16#05#),
      2851 => to_slv(opcode_type, 16#05#),
      2852 => to_slv(opcode_type, 16#0B#),
      2853 => to_slv(opcode_type, 16#09#),
      2854 => to_slv(opcode_type, 16#06#),
      2855 => to_slv(opcode_type, 16#11#),
      2856 => to_slv(opcode_type, 16#F0#),
      2857 => to_slv(opcode_type, 16#07#),
      2858 => to_slv(opcode_type, 16#0F#),
      2859 => to_slv(opcode_type, 16#0F#),
      2860 => to_slv(opcode_type, 16#06#),
      2861 => to_slv(opcode_type, 16#08#),
      2862 => to_slv(opcode_type, 16#09#),
      2863 => to_slv(opcode_type, 16#11#),
      2864 => to_slv(opcode_type, 16#0A#),
      2865 => to_slv(opcode_type, 16#06#),
      2866 => to_slv(opcode_type, 16#0D#),
      2867 => to_slv(opcode_type, 16#0C#),
      2868 => to_slv(opcode_type, 16#07#),
      2869 => to_slv(opcode_type, 16#09#),
      2870 => to_slv(opcode_type, 16#D5#),
      2871 => to_slv(opcode_type, 16#0A#),
      2872 => to_slv(opcode_type, 16#07#),
      2873 => to_slv(opcode_type, 16#0F#),
      2874 => to_slv(opcode_type, 16#1B#),
      2875 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#09#),
      2881 => to_slv(opcode_type, 16#08#),
      2882 => to_slv(opcode_type, 16#07#),
      2883 => to_slv(opcode_type, 16#08#),
      2884 => to_slv(opcode_type, 16#0B#),
      2885 => to_slv(opcode_type, 16#0B#),
      2886 => to_slv(opcode_type, 16#04#),
      2887 => to_slv(opcode_type, 16#10#),
      2888 => to_slv(opcode_type, 16#03#),
      2889 => to_slv(opcode_type, 16#09#),
      2890 => to_slv(opcode_type, 16#50#),
      2891 => to_slv(opcode_type, 16#0D#),
      2892 => to_slv(opcode_type, 16#09#),
      2893 => to_slv(opcode_type, 16#08#),
      2894 => to_slv(opcode_type, 16#08#),
      2895 => to_slv(opcode_type, 16#0F#),
      2896 => to_slv(opcode_type, 16#0C#),
      2897 => to_slv(opcode_type, 16#07#),
      2898 => to_slv(opcode_type, 16#AA#),
      2899 => to_slv(opcode_type, 16#0A#),
      2900 => to_slv(opcode_type, 16#09#),
      2901 => to_slv(opcode_type, 16#06#),
      2902 => to_slv(opcode_type, 16#0C#),
      2903 => to_slv(opcode_type, 16#0E#),
      2904 => to_slv(opcode_type, 16#08#),
      2905 => to_slv(opcode_type, 16#D8#),
      2906 => to_slv(opcode_type, 16#3C#),
      2907 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#09#),
      2913 => to_slv(opcode_type, 16#06#),
      2914 => to_slv(opcode_type, 16#03#),
      2915 => to_slv(opcode_type, 16#07#),
      2916 => to_slv(opcode_type, 16#5F#),
      2917 => to_slv(opcode_type, 16#10#),
      2918 => to_slv(opcode_type, 16#09#),
      2919 => to_slv(opcode_type, 16#09#),
      2920 => to_slv(opcode_type, 16#10#),
      2921 => to_slv(opcode_type, 16#0F#),
      2922 => to_slv(opcode_type, 16#07#),
      2923 => to_slv(opcode_type, 16#11#),
      2924 => to_slv(opcode_type, 16#0A#),
      2925 => to_slv(opcode_type, 16#07#),
      2926 => to_slv(opcode_type, 16#06#),
      2927 => to_slv(opcode_type, 16#08#),
      2928 => to_slv(opcode_type, 16#0E#),
      2929 => to_slv(opcode_type, 16#0F#),
      2930 => to_slv(opcode_type, 16#03#),
      2931 => to_slv(opcode_type, 16#10#),
      2932 => to_slv(opcode_type, 16#06#),
      2933 => to_slv(opcode_type, 16#08#),
      2934 => to_slv(opcode_type, 16#0A#),
      2935 => to_slv(opcode_type, 16#D5#),
      2936 => to_slv(opcode_type, 16#07#),
      2937 => to_slv(opcode_type, 16#0D#),
      2938 => to_slv(opcode_type, 16#0A#),
      2939 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#09#),
      2945 => to_slv(opcode_type, 16#08#),
      2946 => to_slv(opcode_type, 16#02#),
      2947 => to_slv(opcode_type, 16#09#),
      2948 => to_slv(opcode_type, 16#0B#),
      2949 => to_slv(opcode_type, 16#0C#),
      2950 => to_slv(opcode_type, 16#06#),
      2951 => to_slv(opcode_type, 16#08#),
      2952 => to_slv(opcode_type, 16#0D#),
      2953 => to_slv(opcode_type, 16#11#),
      2954 => to_slv(opcode_type, 16#06#),
      2955 => to_slv(opcode_type, 16#0B#),
      2956 => to_slv(opcode_type, 16#0C#),
      2957 => to_slv(opcode_type, 16#08#),
      2958 => to_slv(opcode_type, 16#09#),
      2959 => to_slv(opcode_type, 16#07#),
      2960 => to_slv(opcode_type, 16#F1#),
      2961 => to_slv(opcode_type, 16#D7#),
      2962 => to_slv(opcode_type, 16#05#),
      2963 => to_slv(opcode_type, 16#0E#),
      2964 => to_slv(opcode_type, 16#07#),
      2965 => to_slv(opcode_type, 16#08#),
      2966 => to_slv(opcode_type, 16#0C#),
      2967 => to_slv(opcode_type, 16#0D#),
      2968 => to_slv(opcode_type, 16#08#),
      2969 => to_slv(opcode_type, 16#0F#),
      2970 => to_slv(opcode_type, 16#11#),
      2971 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#06#),
      2977 => to_slv(opcode_type, 16#09#),
      2978 => to_slv(opcode_type, 16#07#),
      2979 => to_slv(opcode_type, 16#04#),
      2980 => to_slv(opcode_type, 16#10#),
      2981 => to_slv(opcode_type, 16#03#),
      2982 => to_slv(opcode_type, 16#0D#),
      2983 => to_slv(opcode_type, 16#09#),
      2984 => to_slv(opcode_type, 16#07#),
      2985 => to_slv(opcode_type, 16#0F#),
      2986 => to_slv(opcode_type, 16#0B#),
      2987 => to_slv(opcode_type, 16#08#),
      2988 => to_slv(opcode_type, 16#0D#),
      2989 => to_slv(opcode_type, 16#BB#),
      2990 => to_slv(opcode_type, 16#08#),
      2991 => to_slv(opcode_type, 16#07#),
      2992 => to_slv(opcode_type, 16#03#),
      2993 => to_slv(opcode_type, 16#0B#),
      2994 => to_slv(opcode_type, 16#03#),
      2995 => to_slv(opcode_type, 16#0E#),
      2996 => to_slv(opcode_type, 16#09#),
      2997 => to_slv(opcode_type, 16#06#),
      2998 => to_slv(opcode_type, 16#0F#),
      2999 => to_slv(opcode_type, 16#0F#),
      3000 => to_slv(opcode_type, 16#09#),
      3001 => to_slv(opcode_type, 16#10#),
      3002 => to_slv(opcode_type, 16#0A#),
      3003 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#07#),
      3009 => to_slv(opcode_type, 16#07#),
      3010 => to_slv(opcode_type, 16#01#),
      3011 => to_slv(opcode_type, 16#03#),
      3012 => to_slv(opcode_type, 16#11#),
      3013 => to_slv(opcode_type, 16#07#),
      3014 => to_slv(opcode_type, 16#07#),
      3015 => to_slv(opcode_type, 16#0E#),
      3016 => to_slv(opcode_type, 16#10#),
      3017 => to_slv(opcode_type, 16#08#),
      3018 => to_slv(opcode_type, 16#0B#),
      3019 => to_slv(opcode_type, 16#0C#),
      3020 => to_slv(opcode_type, 16#06#),
      3021 => to_slv(opcode_type, 16#09#),
      3022 => to_slv(opcode_type, 16#07#),
      3023 => to_slv(opcode_type, 16#0E#),
      3024 => to_slv(opcode_type, 16#11#),
      3025 => to_slv(opcode_type, 16#09#),
      3026 => to_slv(opcode_type, 16#0B#),
      3027 => to_slv(opcode_type, 16#F2#),
      3028 => to_slv(opcode_type, 16#08#),
      3029 => to_slv(opcode_type, 16#06#),
      3030 => to_slv(opcode_type, 16#10#),
      3031 => to_slv(opcode_type, 16#0F#),
      3032 => to_slv(opcode_type, 16#08#),
      3033 => to_slv(opcode_type, 16#0D#),
      3034 => to_slv(opcode_type, 16#10#),
      3035 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#07#),
      3041 => to_slv(opcode_type, 16#09#),
      3042 => to_slv(opcode_type, 16#05#),
      3043 => to_slv(opcode_type, 16#06#),
      3044 => to_slv(opcode_type, 16#0A#),
      3045 => to_slv(opcode_type, 16#0D#),
      3046 => to_slv(opcode_type, 16#09#),
      3047 => to_slv(opcode_type, 16#09#),
      3048 => to_slv(opcode_type, 16#0B#),
      3049 => to_slv(opcode_type, 16#0C#),
      3050 => to_slv(opcode_type, 16#08#),
      3051 => to_slv(opcode_type, 16#0C#),
      3052 => to_slv(opcode_type, 16#0E#),
      3053 => to_slv(opcode_type, 16#07#),
      3054 => to_slv(opcode_type, 16#09#),
      3055 => to_slv(opcode_type, 16#05#),
      3056 => to_slv(opcode_type, 16#4C#),
      3057 => to_slv(opcode_type, 16#07#),
      3058 => to_slv(opcode_type, 16#0C#),
      3059 => to_slv(opcode_type, 16#11#),
      3060 => to_slv(opcode_type, 16#07#),
      3061 => to_slv(opcode_type, 16#07#),
      3062 => to_slv(opcode_type, 16#0B#),
      3063 => to_slv(opcode_type, 16#10#),
      3064 => to_slv(opcode_type, 16#09#),
      3065 => to_slv(opcode_type, 16#0D#),
      3066 => to_slv(opcode_type, 16#0C#),
      3067 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#07#),
      3073 => to_slv(opcode_type, 16#09#),
      3074 => to_slv(opcode_type, 16#05#),
      3075 => to_slv(opcode_type, 16#06#),
      3076 => to_slv(opcode_type, 16#0B#),
      3077 => to_slv(opcode_type, 16#11#),
      3078 => to_slv(opcode_type, 16#08#),
      3079 => to_slv(opcode_type, 16#06#),
      3080 => to_slv(opcode_type, 16#0F#),
      3081 => to_slv(opcode_type, 16#0D#),
      3082 => to_slv(opcode_type, 16#09#),
      3083 => to_slv(opcode_type, 16#10#),
      3084 => to_slv(opcode_type, 16#10#),
      3085 => to_slv(opcode_type, 16#08#),
      3086 => to_slv(opcode_type, 16#08#),
      3087 => to_slv(opcode_type, 16#02#),
      3088 => to_slv(opcode_type, 16#10#),
      3089 => to_slv(opcode_type, 16#09#),
      3090 => to_slv(opcode_type, 16#0D#),
      3091 => to_slv(opcode_type, 16#11#),
      3092 => to_slv(opcode_type, 16#06#),
      3093 => to_slv(opcode_type, 16#08#),
      3094 => to_slv(opcode_type, 16#11#),
      3095 => to_slv(opcode_type, 16#0E#),
      3096 => to_slv(opcode_type, 16#07#),
      3097 => to_slv(opcode_type, 16#0A#),
      3098 => to_slv(opcode_type, 16#0D#),
      3099 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#06#),
      3105 => to_slv(opcode_type, 16#09#),
      3106 => to_slv(opcode_type, 16#05#),
      3107 => to_slv(opcode_type, 16#08#),
      3108 => to_slv(opcode_type, 16#0D#),
      3109 => to_slv(opcode_type, 16#6D#),
      3110 => to_slv(opcode_type, 16#09#),
      3111 => to_slv(opcode_type, 16#04#),
      3112 => to_slv(opcode_type, 16#10#),
      3113 => to_slv(opcode_type, 16#07#),
      3114 => to_slv(opcode_type, 16#10#),
      3115 => to_slv(opcode_type, 16#AB#),
      3116 => to_slv(opcode_type, 16#06#),
      3117 => to_slv(opcode_type, 16#08#),
      3118 => to_slv(opcode_type, 16#06#),
      3119 => to_slv(opcode_type, 16#0D#),
      3120 => to_slv(opcode_type, 16#10#),
      3121 => to_slv(opcode_type, 16#09#),
      3122 => to_slv(opcode_type, 16#0B#),
      3123 => to_slv(opcode_type, 16#0B#),
      3124 => to_slv(opcode_type, 16#08#),
      3125 => to_slv(opcode_type, 16#09#),
      3126 => to_slv(opcode_type, 16#0A#),
      3127 => to_slv(opcode_type, 16#0D#),
      3128 => to_slv(opcode_type, 16#07#),
      3129 => to_slv(opcode_type, 16#0A#),
      3130 => to_slv(opcode_type, 16#82#),
      3131 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#06#),
      3137 => to_slv(opcode_type, 16#06#),
      3138 => to_slv(opcode_type, 16#03#),
      3139 => to_slv(opcode_type, 16#05#),
      3140 => to_slv(opcode_type, 16#0A#),
      3141 => to_slv(opcode_type, 16#08#),
      3142 => to_slv(opcode_type, 16#08#),
      3143 => to_slv(opcode_type, 16#11#),
      3144 => to_slv(opcode_type, 16#0B#),
      3145 => to_slv(opcode_type, 16#09#),
      3146 => to_slv(opcode_type, 16#11#),
      3147 => to_slv(opcode_type, 16#11#),
      3148 => to_slv(opcode_type, 16#09#),
      3149 => to_slv(opcode_type, 16#09#),
      3150 => to_slv(opcode_type, 16#07#),
      3151 => to_slv(opcode_type, 16#0F#),
      3152 => to_slv(opcode_type, 16#0A#),
      3153 => to_slv(opcode_type, 16#09#),
      3154 => to_slv(opcode_type, 16#11#),
      3155 => to_slv(opcode_type, 16#0C#),
      3156 => to_slv(opcode_type, 16#08#),
      3157 => to_slv(opcode_type, 16#06#),
      3158 => to_slv(opcode_type, 16#0F#),
      3159 => to_slv(opcode_type, 16#11#),
      3160 => to_slv(opcode_type, 16#09#),
      3161 => to_slv(opcode_type, 16#0D#),
      3162 => to_slv(opcode_type, 16#0A#),
      3163 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#07#),
      3169 => to_slv(opcode_type, 16#08#),
      3170 => to_slv(opcode_type, 16#03#),
      3171 => to_slv(opcode_type, 16#07#),
      3172 => to_slv(opcode_type, 16#0B#),
      3173 => to_slv(opcode_type, 16#0D#),
      3174 => to_slv(opcode_type, 16#07#),
      3175 => to_slv(opcode_type, 16#09#),
      3176 => to_slv(opcode_type, 16#0D#),
      3177 => to_slv(opcode_type, 16#EF#),
      3178 => to_slv(opcode_type, 16#03#),
      3179 => to_slv(opcode_type, 16#0A#),
      3180 => to_slv(opcode_type, 16#07#),
      3181 => to_slv(opcode_type, 16#06#),
      3182 => to_slv(opcode_type, 16#09#),
      3183 => to_slv(opcode_type, 16#0F#),
      3184 => to_slv(opcode_type, 16#10#),
      3185 => to_slv(opcode_type, 16#06#),
      3186 => to_slv(opcode_type, 16#60#),
      3187 => to_slv(opcode_type, 16#11#),
      3188 => to_slv(opcode_type, 16#08#),
      3189 => to_slv(opcode_type, 16#09#),
      3190 => to_slv(opcode_type, 16#0D#),
      3191 => to_slv(opcode_type, 16#0C#),
      3192 => to_slv(opcode_type, 16#09#),
      3193 => to_slv(opcode_type, 16#11#),
      3194 => to_slv(opcode_type, 16#10#),
      3195 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#09#),
      3201 => to_slv(opcode_type, 16#08#),
      3202 => to_slv(opcode_type, 16#06#),
      3203 => to_slv(opcode_type, 16#09#),
      3204 => to_slv(opcode_type, 16#11#),
      3205 => to_slv(opcode_type, 16#0F#),
      3206 => to_slv(opcode_type, 16#05#),
      3207 => to_slv(opcode_type, 16#91#),
      3208 => to_slv(opcode_type, 16#01#),
      3209 => to_slv(opcode_type, 16#07#),
      3210 => to_slv(opcode_type, 16#C5#),
      3211 => to_slv(opcode_type, 16#0F#),
      3212 => to_slv(opcode_type, 16#06#),
      3213 => to_slv(opcode_type, 16#09#),
      3214 => to_slv(opcode_type, 16#08#),
      3215 => to_slv(opcode_type, 16#0E#),
      3216 => to_slv(opcode_type, 16#0B#),
      3217 => to_slv(opcode_type, 16#06#),
      3218 => to_slv(opcode_type, 16#0A#),
      3219 => to_slv(opcode_type, 16#0B#),
      3220 => to_slv(opcode_type, 16#08#),
      3221 => to_slv(opcode_type, 16#08#),
      3222 => to_slv(opcode_type, 16#10#),
      3223 => to_slv(opcode_type, 16#0B#),
      3224 => to_slv(opcode_type, 16#08#),
      3225 => to_slv(opcode_type, 16#0C#),
      3226 => to_slv(opcode_type, 16#89#),
      3227 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#07#),
      3234 => to_slv(opcode_type, 16#05#),
      3235 => to_slv(opcode_type, 16#03#),
      3236 => to_slv(opcode_type, 16#0B#),
      3237 => to_slv(opcode_type, 16#06#),
      3238 => to_slv(opcode_type, 16#06#),
      3239 => to_slv(opcode_type, 16#0E#),
      3240 => to_slv(opcode_type, 16#11#),
      3241 => to_slv(opcode_type, 16#06#),
      3242 => to_slv(opcode_type, 16#0D#),
      3243 => to_slv(opcode_type, 16#11#),
      3244 => to_slv(opcode_type, 16#09#),
      3245 => to_slv(opcode_type, 16#09#),
      3246 => to_slv(opcode_type, 16#08#),
      3247 => to_slv(opcode_type, 16#0A#),
      3248 => to_slv(opcode_type, 16#10#),
      3249 => to_slv(opcode_type, 16#08#),
      3250 => to_slv(opcode_type, 16#11#),
      3251 => to_slv(opcode_type, 16#0B#),
      3252 => to_slv(opcode_type, 16#07#),
      3253 => to_slv(opcode_type, 16#08#),
      3254 => to_slv(opcode_type, 16#0B#),
      3255 => to_slv(opcode_type, 16#0F#),
      3256 => to_slv(opcode_type, 16#09#),
      3257 => to_slv(opcode_type, 16#0D#),
      3258 => to_slv(opcode_type, 16#40#),
      3259 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#09#),
      3265 => to_slv(opcode_type, 16#06#),
      3266 => to_slv(opcode_type, 16#02#),
      3267 => to_slv(opcode_type, 16#08#),
      3268 => to_slv(opcode_type, 16#11#),
      3269 => to_slv(opcode_type, 16#10#),
      3270 => to_slv(opcode_type, 16#07#),
      3271 => to_slv(opcode_type, 16#06#),
      3272 => to_slv(opcode_type, 16#31#),
      3273 => to_slv(opcode_type, 16#0C#),
      3274 => to_slv(opcode_type, 16#03#),
      3275 => to_slv(opcode_type, 16#73#),
      3276 => to_slv(opcode_type, 16#08#),
      3277 => to_slv(opcode_type, 16#09#),
      3278 => to_slv(opcode_type, 16#07#),
      3279 => to_slv(opcode_type, 16#0E#),
      3280 => to_slv(opcode_type, 16#11#),
      3281 => to_slv(opcode_type, 16#09#),
      3282 => to_slv(opcode_type, 16#11#),
      3283 => to_slv(opcode_type, 16#0F#),
      3284 => to_slv(opcode_type, 16#09#),
      3285 => to_slv(opcode_type, 16#06#),
      3286 => to_slv(opcode_type, 16#BD#),
      3287 => to_slv(opcode_type, 16#10#),
      3288 => to_slv(opcode_type, 16#09#),
      3289 => to_slv(opcode_type, 16#3F#),
      3290 => to_slv(opcode_type, 16#0D#),
      3291 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#09#),
      3297 => to_slv(opcode_type, 16#07#),
      3298 => to_slv(opcode_type, 16#08#),
      3299 => to_slv(opcode_type, 16#06#),
      3300 => to_slv(opcode_type, 16#CD#),
      3301 => to_slv(opcode_type, 16#0E#),
      3302 => to_slv(opcode_type, 16#05#),
      3303 => to_slv(opcode_type, 16#0E#),
      3304 => to_slv(opcode_type, 16#03#),
      3305 => to_slv(opcode_type, 16#09#),
      3306 => to_slv(opcode_type, 16#0F#),
      3307 => to_slv(opcode_type, 16#0A#),
      3308 => to_slv(opcode_type, 16#09#),
      3309 => to_slv(opcode_type, 16#06#),
      3310 => to_slv(opcode_type, 16#09#),
      3311 => to_slv(opcode_type, 16#E5#),
      3312 => to_slv(opcode_type, 16#11#),
      3313 => to_slv(opcode_type, 16#07#),
      3314 => to_slv(opcode_type, 16#11#),
      3315 => to_slv(opcode_type, 16#0D#),
      3316 => to_slv(opcode_type, 16#06#),
      3317 => to_slv(opcode_type, 16#08#),
      3318 => to_slv(opcode_type, 16#0E#),
      3319 => to_slv(opcode_type, 16#0B#),
      3320 => to_slv(opcode_type, 16#07#),
      3321 => to_slv(opcode_type, 16#0C#),
      3322 => to_slv(opcode_type, 16#11#),
      3323 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#09#),
      3329 => to_slv(opcode_type, 16#08#),
      3330 => to_slv(opcode_type, 16#02#),
      3331 => to_slv(opcode_type, 16#07#),
      3332 => to_slv(opcode_type, 16#0E#),
      3333 => to_slv(opcode_type, 16#10#),
      3334 => to_slv(opcode_type, 16#07#),
      3335 => to_slv(opcode_type, 16#05#),
      3336 => to_slv(opcode_type, 16#0D#),
      3337 => to_slv(opcode_type, 16#06#),
      3338 => to_slv(opcode_type, 16#0E#),
      3339 => to_slv(opcode_type, 16#0E#),
      3340 => to_slv(opcode_type, 16#06#),
      3341 => to_slv(opcode_type, 16#08#),
      3342 => to_slv(opcode_type, 16#09#),
      3343 => to_slv(opcode_type, 16#0F#),
      3344 => to_slv(opcode_type, 16#0E#),
      3345 => to_slv(opcode_type, 16#07#),
      3346 => to_slv(opcode_type, 16#2B#),
      3347 => to_slv(opcode_type, 16#0C#),
      3348 => to_slv(opcode_type, 16#09#),
      3349 => to_slv(opcode_type, 16#09#),
      3350 => to_slv(opcode_type, 16#11#),
      3351 => to_slv(opcode_type, 16#46#),
      3352 => to_slv(opcode_type, 16#09#),
      3353 => to_slv(opcode_type, 16#0B#),
      3354 => to_slv(opcode_type, 16#0E#),
      3355 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#08#),
      3361 => to_slv(opcode_type, 16#08#),
      3362 => to_slv(opcode_type, 16#08#),
      3363 => to_slv(opcode_type, 16#07#),
      3364 => to_slv(opcode_type, 16#0B#),
      3365 => to_slv(opcode_type, 16#0E#),
      3366 => to_slv(opcode_type, 16#08#),
      3367 => to_slv(opcode_type, 16#0E#),
      3368 => to_slv(opcode_type, 16#0D#),
      3369 => to_slv(opcode_type, 16#04#),
      3370 => to_slv(opcode_type, 16#07#),
      3371 => to_slv(opcode_type, 16#0E#),
      3372 => to_slv(opcode_type, 16#10#),
      3373 => to_slv(opcode_type, 16#06#),
      3374 => to_slv(opcode_type, 16#07#),
      3375 => to_slv(opcode_type, 16#02#),
      3376 => to_slv(opcode_type, 16#0B#),
      3377 => to_slv(opcode_type, 16#08#),
      3378 => to_slv(opcode_type, 16#0D#),
      3379 => to_slv(opcode_type, 16#0E#),
      3380 => to_slv(opcode_type, 16#07#),
      3381 => to_slv(opcode_type, 16#09#),
      3382 => to_slv(opcode_type, 16#11#),
      3383 => to_slv(opcode_type, 16#0E#),
      3384 => to_slv(opcode_type, 16#06#),
      3385 => to_slv(opcode_type, 16#11#),
      3386 => to_slv(opcode_type, 16#CB#),
      3387 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#08#),
      3393 => to_slv(opcode_type, 16#07#),
      3394 => to_slv(opcode_type, 16#02#),
      3395 => to_slv(opcode_type, 16#09#),
      3396 => to_slv(opcode_type, 16#0E#),
      3397 => to_slv(opcode_type, 16#0D#),
      3398 => to_slv(opcode_type, 16#06#),
      3399 => to_slv(opcode_type, 16#05#),
      3400 => to_slv(opcode_type, 16#0B#),
      3401 => to_slv(opcode_type, 16#06#),
      3402 => to_slv(opcode_type, 16#11#),
      3403 => to_slv(opcode_type, 16#82#),
      3404 => to_slv(opcode_type, 16#07#),
      3405 => to_slv(opcode_type, 16#09#),
      3406 => to_slv(opcode_type, 16#09#),
      3407 => to_slv(opcode_type, 16#0E#),
      3408 => to_slv(opcode_type, 16#0A#),
      3409 => to_slv(opcode_type, 16#07#),
      3410 => to_slv(opcode_type, 16#10#),
      3411 => to_slv(opcode_type, 16#0F#),
      3412 => to_slv(opcode_type, 16#07#),
      3413 => to_slv(opcode_type, 16#06#),
      3414 => to_slv(opcode_type, 16#0A#),
      3415 => to_slv(opcode_type, 16#0E#),
      3416 => to_slv(opcode_type, 16#08#),
      3417 => to_slv(opcode_type, 16#0C#),
      3418 => to_slv(opcode_type, 16#0A#),
      3419 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#09#),
      3425 => to_slv(opcode_type, 16#09#),
      3426 => to_slv(opcode_type, 16#04#),
      3427 => to_slv(opcode_type, 16#02#),
      3428 => to_slv(opcode_type, 16#34#),
      3429 => to_slv(opcode_type, 16#06#),
      3430 => to_slv(opcode_type, 16#09#),
      3431 => to_slv(opcode_type, 16#0B#),
      3432 => to_slv(opcode_type, 16#0E#),
      3433 => to_slv(opcode_type, 16#07#),
      3434 => to_slv(opcode_type, 16#0E#),
      3435 => to_slv(opcode_type, 16#0F#),
      3436 => to_slv(opcode_type, 16#06#),
      3437 => to_slv(opcode_type, 16#08#),
      3438 => to_slv(opcode_type, 16#08#),
      3439 => to_slv(opcode_type, 16#0E#),
      3440 => to_slv(opcode_type, 16#11#),
      3441 => to_slv(opcode_type, 16#08#),
      3442 => to_slv(opcode_type, 16#0F#),
      3443 => to_slv(opcode_type, 16#0C#),
      3444 => to_slv(opcode_type, 16#06#),
      3445 => to_slv(opcode_type, 16#09#),
      3446 => to_slv(opcode_type, 16#11#),
      3447 => to_slv(opcode_type, 16#0E#),
      3448 => to_slv(opcode_type, 16#09#),
      3449 => to_slv(opcode_type, 16#0F#),
      3450 => to_slv(opcode_type, 16#86#),
      3451 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#08#),
      3457 => to_slv(opcode_type, 16#09#),
      3458 => to_slv(opcode_type, 16#04#),
      3459 => to_slv(opcode_type, 16#07#),
      3460 => to_slv(opcode_type, 16#0C#),
      3461 => to_slv(opcode_type, 16#0F#),
      3462 => to_slv(opcode_type, 16#08#),
      3463 => to_slv(opcode_type, 16#05#),
      3464 => to_slv(opcode_type, 16#BD#),
      3465 => to_slv(opcode_type, 16#06#),
      3466 => to_slv(opcode_type, 16#40#),
      3467 => to_slv(opcode_type, 16#0C#),
      3468 => to_slv(opcode_type, 16#09#),
      3469 => to_slv(opcode_type, 16#07#),
      3470 => to_slv(opcode_type, 16#08#),
      3471 => to_slv(opcode_type, 16#0F#),
      3472 => to_slv(opcode_type, 16#DC#),
      3473 => to_slv(opcode_type, 16#07#),
      3474 => to_slv(opcode_type, 16#0B#),
      3475 => to_slv(opcode_type, 16#0A#),
      3476 => to_slv(opcode_type, 16#08#),
      3477 => to_slv(opcode_type, 16#06#),
      3478 => to_slv(opcode_type, 16#0A#),
      3479 => to_slv(opcode_type, 16#11#),
      3480 => to_slv(opcode_type, 16#08#),
      3481 => to_slv(opcode_type, 16#11#),
      3482 => to_slv(opcode_type, 16#10#),
      3483 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#07#),
      3489 => to_slv(opcode_type, 16#08#),
      3490 => to_slv(opcode_type, 16#07#),
      3491 => to_slv(opcode_type, 16#02#),
      3492 => to_slv(opcode_type, 16#0C#),
      3493 => to_slv(opcode_type, 16#04#),
      3494 => to_slv(opcode_type, 16#0E#),
      3495 => to_slv(opcode_type, 16#07#),
      3496 => to_slv(opcode_type, 16#03#),
      3497 => to_slv(opcode_type, 16#0E#),
      3498 => to_slv(opcode_type, 16#03#),
      3499 => to_slv(opcode_type, 16#0F#),
      3500 => to_slv(opcode_type, 16#08#),
      3501 => to_slv(opcode_type, 16#06#),
      3502 => to_slv(opcode_type, 16#06#),
      3503 => to_slv(opcode_type, 16#0A#),
      3504 => to_slv(opcode_type, 16#0E#),
      3505 => to_slv(opcode_type, 16#08#),
      3506 => to_slv(opcode_type, 16#0B#),
      3507 => to_slv(opcode_type, 16#FC#),
      3508 => to_slv(opcode_type, 16#06#),
      3509 => to_slv(opcode_type, 16#06#),
      3510 => to_slv(opcode_type, 16#0A#),
      3511 => to_slv(opcode_type, 16#11#),
      3512 => to_slv(opcode_type, 16#07#),
      3513 => to_slv(opcode_type, 16#0A#),
      3514 => to_slv(opcode_type, 16#0C#),
      3515 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#09#),
      3521 => to_slv(opcode_type, 16#08#),
      3522 => to_slv(opcode_type, 16#01#),
      3523 => to_slv(opcode_type, 16#07#),
      3524 => to_slv(opcode_type, 16#11#),
      3525 => to_slv(opcode_type, 16#0E#),
      3526 => to_slv(opcode_type, 16#08#),
      3527 => to_slv(opcode_type, 16#04#),
      3528 => to_slv(opcode_type, 16#0A#),
      3529 => to_slv(opcode_type, 16#09#),
      3530 => to_slv(opcode_type, 16#0E#),
      3531 => to_slv(opcode_type, 16#0C#),
      3532 => to_slv(opcode_type, 16#08#),
      3533 => to_slv(opcode_type, 16#06#),
      3534 => to_slv(opcode_type, 16#07#),
      3535 => to_slv(opcode_type, 16#0E#),
      3536 => to_slv(opcode_type, 16#0C#),
      3537 => to_slv(opcode_type, 16#09#),
      3538 => to_slv(opcode_type, 16#0E#),
      3539 => to_slv(opcode_type, 16#11#),
      3540 => to_slv(opcode_type, 16#07#),
      3541 => to_slv(opcode_type, 16#07#),
      3542 => to_slv(opcode_type, 16#0E#),
      3543 => to_slv(opcode_type, 16#10#),
      3544 => to_slv(opcode_type, 16#07#),
      3545 => to_slv(opcode_type, 16#0E#),
      3546 => to_slv(opcode_type, 16#0F#),
      3547 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#06#),
      3553 => to_slv(opcode_type, 16#07#),
      3554 => to_slv(opcode_type, 16#07#),
      3555 => to_slv(opcode_type, 16#06#),
      3556 => to_slv(opcode_type, 16#10#),
      3557 => to_slv(opcode_type, 16#0E#),
      3558 => to_slv(opcode_type, 16#05#),
      3559 => to_slv(opcode_type, 16#10#),
      3560 => to_slv(opcode_type, 16#03#),
      3561 => to_slv(opcode_type, 16#08#),
      3562 => to_slv(opcode_type, 16#74#),
      3563 => to_slv(opcode_type, 16#0E#),
      3564 => to_slv(opcode_type, 16#09#),
      3565 => to_slv(opcode_type, 16#07#),
      3566 => to_slv(opcode_type, 16#06#),
      3567 => to_slv(opcode_type, 16#0C#),
      3568 => to_slv(opcode_type, 16#0C#),
      3569 => to_slv(opcode_type, 16#09#),
      3570 => to_slv(opcode_type, 16#0D#),
      3571 => to_slv(opcode_type, 16#0F#),
      3572 => to_slv(opcode_type, 16#06#),
      3573 => to_slv(opcode_type, 16#07#),
      3574 => to_slv(opcode_type, 16#0B#),
      3575 => to_slv(opcode_type, 16#0B#),
      3576 => to_slv(opcode_type, 16#07#),
      3577 => to_slv(opcode_type, 16#0D#),
      3578 => to_slv(opcode_type, 16#0B#),
      3579 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#09#),
      3585 => to_slv(opcode_type, 16#07#),
      3586 => to_slv(opcode_type, 16#07#),
      3587 => to_slv(opcode_type, 16#07#),
      3588 => to_slv(opcode_type, 16#0E#),
      3589 => to_slv(opcode_type, 16#0A#),
      3590 => to_slv(opcode_type, 16#05#),
      3591 => to_slv(opcode_type, 16#10#),
      3592 => to_slv(opcode_type, 16#08#),
      3593 => to_slv(opcode_type, 16#07#),
      3594 => to_slv(opcode_type, 16#0B#),
      3595 => to_slv(opcode_type, 16#0B#),
      3596 => to_slv(opcode_type, 16#06#),
      3597 => to_slv(opcode_type, 16#11#),
      3598 => to_slv(opcode_type, 16#0A#),
      3599 => to_slv(opcode_type, 16#08#),
      3600 => to_slv(opcode_type, 16#07#),
      3601 => to_slv(opcode_type, 16#08#),
      3602 => to_slv(opcode_type, 16#0B#),
      3603 => to_slv(opcode_type, 16#0A#),
      3604 => to_slv(opcode_type, 16#04#),
      3605 => to_slv(opcode_type, 16#0F#),
      3606 => to_slv(opcode_type, 16#09#),
      3607 => to_slv(opcode_type, 16#02#),
      3608 => to_slv(opcode_type, 16#0E#),
      3609 => to_slv(opcode_type, 16#02#),
      3610 => to_slv(opcode_type, 16#5D#),
      3611 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#07#),
      3617 => to_slv(opcode_type, 16#09#),
      3618 => to_slv(opcode_type, 16#04#),
      3619 => to_slv(opcode_type, 16#08#),
      3620 => to_slv(opcode_type, 16#0E#),
      3621 => to_slv(opcode_type, 16#10#),
      3622 => to_slv(opcode_type, 16#09#),
      3623 => to_slv(opcode_type, 16#01#),
      3624 => to_slv(opcode_type, 16#0F#),
      3625 => to_slv(opcode_type, 16#06#),
      3626 => to_slv(opcode_type, 16#0F#),
      3627 => to_slv(opcode_type, 16#0F#),
      3628 => to_slv(opcode_type, 16#08#),
      3629 => to_slv(opcode_type, 16#09#),
      3630 => to_slv(opcode_type, 16#06#),
      3631 => to_slv(opcode_type, 16#0D#),
      3632 => to_slv(opcode_type, 16#0E#),
      3633 => to_slv(opcode_type, 16#07#),
      3634 => to_slv(opcode_type, 16#0B#),
      3635 => to_slv(opcode_type, 16#0D#),
      3636 => to_slv(opcode_type, 16#07#),
      3637 => to_slv(opcode_type, 16#06#),
      3638 => to_slv(opcode_type, 16#0A#),
      3639 => to_slv(opcode_type, 16#0A#),
      3640 => to_slv(opcode_type, 16#07#),
      3641 => to_slv(opcode_type, 16#11#),
      3642 => to_slv(opcode_type, 16#0C#),
      3643 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#07#),
      3649 => to_slv(opcode_type, 16#09#),
      3650 => to_slv(opcode_type, 16#05#),
      3651 => to_slv(opcode_type, 16#05#),
      3652 => to_slv(opcode_type, 16#0F#),
      3653 => to_slv(opcode_type, 16#06#),
      3654 => to_slv(opcode_type, 16#07#),
      3655 => to_slv(opcode_type, 16#0F#),
      3656 => to_slv(opcode_type, 16#11#),
      3657 => to_slv(opcode_type, 16#09#),
      3658 => to_slv(opcode_type, 16#0C#),
      3659 => to_slv(opcode_type, 16#37#),
      3660 => to_slv(opcode_type, 16#09#),
      3661 => to_slv(opcode_type, 16#09#),
      3662 => to_slv(opcode_type, 16#09#),
      3663 => to_slv(opcode_type, 16#10#),
      3664 => to_slv(opcode_type, 16#0B#),
      3665 => to_slv(opcode_type, 16#08#),
      3666 => to_slv(opcode_type, 16#0D#),
      3667 => to_slv(opcode_type, 16#0F#),
      3668 => to_slv(opcode_type, 16#06#),
      3669 => to_slv(opcode_type, 16#08#),
      3670 => to_slv(opcode_type, 16#45#),
      3671 => to_slv(opcode_type, 16#0B#),
      3672 => to_slv(opcode_type, 16#09#),
      3673 => to_slv(opcode_type, 16#0C#),
      3674 => to_slv(opcode_type, 16#FB#),
      3675 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#06#),
      3681 => to_slv(opcode_type, 16#09#),
      3682 => to_slv(opcode_type, 16#08#),
      3683 => to_slv(opcode_type, 16#07#),
      3684 => to_slv(opcode_type, 16#0C#),
      3685 => to_slv(opcode_type, 16#57#),
      3686 => to_slv(opcode_type, 16#02#),
      3687 => to_slv(opcode_type, 16#10#),
      3688 => to_slv(opcode_type, 16#01#),
      3689 => to_slv(opcode_type, 16#06#),
      3690 => to_slv(opcode_type, 16#11#),
      3691 => to_slv(opcode_type, 16#0B#),
      3692 => to_slv(opcode_type, 16#09#),
      3693 => to_slv(opcode_type, 16#08#),
      3694 => to_slv(opcode_type, 16#07#),
      3695 => to_slv(opcode_type, 16#0A#),
      3696 => to_slv(opcode_type, 16#0E#),
      3697 => to_slv(opcode_type, 16#07#),
      3698 => to_slv(opcode_type, 16#0C#),
      3699 => to_slv(opcode_type, 16#0E#),
      3700 => to_slv(opcode_type, 16#06#),
      3701 => to_slv(opcode_type, 16#08#),
      3702 => to_slv(opcode_type, 16#0A#),
      3703 => to_slv(opcode_type, 16#10#),
      3704 => to_slv(opcode_type, 16#08#),
      3705 => to_slv(opcode_type, 16#0A#),
      3706 => to_slv(opcode_type, 16#0E#),
      3707 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#08#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#09#),
      3715 => to_slv(opcode_type, 16#05#),
      3716 => to_slv(opcode_type, 16#0F#),
      3717 => to_slv(opcode_type, 16#03#),
      3718 => to_slv(opcode_type, 16#0B#),
      3719 => to_slv(opcode_type, 16#07#),
      3720 => to_slv(opcode_type, 16#07#),
      3721 => to_slv(opcode_type, 16#0B#),
      3722 => to_slv(opcode_type, 16#0D#),
      3723 => to_slv(opcode_type, 16#01#),
      3724 => to_slv(opcode_type, 16#0F#),
      3725 => to_slv(opcode_type, 16#08#),
      3726 => to_slv(opcode_type, 16#06#),
      3727 => to_slv(opcode_type, 16#07#),
      3728 => to_slv(opcode_type, 16#0C#),
      3729 => to_slv(opcode_type, 16#0F#),
      3730 => to_slv(opcode_type, 16#06#),
      3731 => to_slv(opcode_type, 16#11#),
      3732 => to_slv(opcode_type, 16#0C#),
      3733 => to_slv(opcode_type, 16#06#),
      3734 => to_slv(opcode_type, 16#07#),
      3735 => to_slv(opcode_type, 16#10#),
      3736 => to_slv(opcode_type, 16#0C#),
      3737 => to_slv(opcode_type, 16#02#),
      3738 => to_slv(opcode_type, 16#6A#),
      3739 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#07#),
      3745 => to_slv(opcode_type, 16#06#),
      3746 => to_slv(opcode_type, 16#09#),
      3747 => to_slv(opcode_type, 16#05#),
      3748 => to_slv(opcode_type, 16#0C#),
      3749 => to_slv(opcode_type, 16#07#),
      3750 => to_slv(opcode_type, 16#0C#),
      3751 => to_slv(opcode_type, 16#10#),
      3752 => to_slv(opcode_type, 16#01#),
      3753 => to_slv(opcode_type, 16#06#),
      3754 => to_slv(opcode_type, 16#10#),
      3755 => to_slv(opcode_type, 16#0A#),
      3756 => to_slv(opcode_type, 16#06#),
      3757 => to_slv(opcode_type, 16#08#),
      3758 => to_slv(opcode_type, 16#06#),
      3759 => to_slv(opcode_type, 16#0E#),
      3760 => to_slv(opcode_type, 16#0D#),
      3761 => to_slv(opcode_type, 16#06#),
      3762 => to_slv(opcode_type, 16#10#),
      3763 => to_slv(opcode_type, 16#0C#),
      3764 => to_slv(opcode_type, 16#09#),
      3765 => to_slv(opcode_type, 16#09#),
      3766 => to_slv(opcode_type, 16#10#),
      3767 => to_slv(opcode_type, 16#11#),
      3768 => to_slv(opcode_type, 16#07#),
      3769 => to_slv(opcode_type, 16#0B#),
      3770 => to_slv(opcode_type, 16#10#),
      3771 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#08#),
      3777 => to_slv(opcode_type, 16#09#),
      3778 => to_slv(opcode_type, 16#05#),
      3779 => to_slv(opcode_type, 16#09#),
      3780 => to_slv(opcode_type, 16#0E#),
      3781 => to_slv(opcode_type, 16#0A#),
      3782 => to_slv(opcode_type, 16#09#),
      3783 => to_slv(opcode_type, 16#02#),
      3784 => to_slv(opcode_type, 16#0C#),
      3785 => to_slv(opcode_type, 16#08#),
      3786 => to_slv(opcode_type, 16#0C#),
      3787 => to_slv(opcode_type, 16#0D#),
      3788 => to_slv(opcode_type, 16#09#),
      3789 => to_slv(opcode_type, 16#08#),
      3790 => to_slv(opcode_type, 16#08#),
      3791 => to_slv(opcode_type, 16#10#),
      3792 => to_slv(opcode_type, 16#0E#),
      3793 => to_slv(opcode_type, 16#07#),
      3794 => to_slv(opcode_type, 16#10#),
      3795 => to_slv(opcode_type, 16#0E#),
      3796 => to_slv(opcode_type, 16#09#),
      3797 => to_slv(opcode_type, 16#08#),
      3798 => to_slv(opcode_type, 16#0F#),
      3799 => to_slv(opcode_type, 16#0E#),
      3800 => to_slv(opcode_type, 16#07#),
      3801 => to_slv(opcode_type, 16#0C#),
      3802 => to_slv(opcode_type, 16#10#),
      3803 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#08#),
      3809 => to_slv(opcode_type, 16#09#),
      3810 => to_slv(opcode_type, 16#08#),
      3811 => to_slv(opcode_type, 16#06#),
      3812 => to_slv(opcode_type, 16#10#),
      3813 => to_slv(opcode_type, 16#0B#),
      3814 => to_slv(opcode_type, 16#02#),
      3815 => to_slv(opcode_type, 16#0C#),
      3816 => to_slv(opcode_type, 16#05#),
      3817 => to_slv(opcode_type, 16#08#),
      3818 => to_slv(opcode_type, 16#0C#),
      3819 => to_slv(opcode_type, 16#11#),
      3820 => to_slv(opcode_type, 16#09#),
      3821 => to_slv(opcode_type, 16#06#),
      3822 => to_slv(opcode_type, 16#06#),
      3823 => to_slv(opcode_type, 16#0A#),
      3824 => to_slv(opcode_type, 16#0A#),
      3825 => to_slv(opcode_type, 16#06#),
      3826 => to_slv(opcode_type, 16#0A#),
      3827 => to_slv(opcode_type, 16#0C#),
      3828 => to_slv(opcode_type, 16#07#),
      3829 => to_slv(opcode_type, 16#07#),
      3830 => to_slv(opcode_type, 16#0E#),
      3831 => to_slv(opcode_type, 16#10#),
      3832 => to_slv(opcode_type, 16#07#),
      3833 => to_slv(opcode_type, 16#33#),
      3834 => to_slv(opcode_type, 16#A5#),
      3835 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#08#),
      3841 => to_slv(opcode_type, 16#06#),
      3842 => to_slv(opcode_type, 16#08#),
      3843 => to_slv(opcode_type, 16#03#),
      3844 => to_slv(opcode_type, 16#10#),
      3845 => to_slv(opcode_type, 16#02#),
      3846 => to_slv(opcode_type, 16#11#),
      3847 => to_slv(opcode_type, 16#08#),
      3848 => to_slv(opcode_type, 16#03#),
      3849 => to_slv(opcode_type, 16#10#),
      3850 => to_slv(opcode_type, 16#08#),
      3851 => to_slv(opcode_type, 16#0E#),
      3852 => to_slv(opcode_type, 16#11#),
      3853 => to_slv(opcode_type, 16#09#),
      3854 => to_slv(opcode_type, 16#08#),
      3855 => to_slv(opcode_type, 16#01#),
      3856 => to_slv(opcode_type, 16#0C#),
      3857 => to_slv(opcode_type, 16#09#),
      3858 => to_slv(opcode_type, 16#0B#),
      3859 => to_slv(opcode_type, 16#10#),
      3860 => to_slv(opcode_type, 16#06#),
      3861 => to_slv(opcode_type, 16#08#),
      3862 => to_slv(opcode_type, 16#8C#),
      3863 => to_slv(opcode_type, 16#11#),
      3864 => to_slv(opcode_type, 16#07#),
      3865 => to_slv(opcode_type, 16#0C#),
      3866 => to_slv(opcode_type, 16#0B#),
      3867 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#09#),
      3873 => to_slv(opcode_type, 16#07#),
      3874 => to_slv(opcode_type, 16#02#),
      3875 => to_slv(opcode_type, 16#09#),
      3876 => to_slv(opcode_type, 16#0B#),
      3877 => to_slv(opcode_type, 16#0D#),
      3878 => to_slv(opcode_type, 16#08#),
      3879 => to_slv(opcode_type, 16#01#),
      3880 => to_slv(opcode_type, 16#0E#),
      3881 => to_slv(opcode_type, 16#08#),
      3882 => to_slv(opcode_type, 16#10#),
      3883 => to_slv(opcode_type, 16#11#),
      3884 => to_slv(opcode_type, 16#09#),
      3885 => to_slv(opcode_type, 16#06#),
      3886 => to_slv(opcode_type, 16#07#),
      3887 => to_slv(opcode_type, 16#0B#),
      3888 => to_slv(opcode_type, 16#3C#),
      3889 => to_slv(opcode_type, 16#09#),
      3890 => to_slv(opcode_type, 16#10#),
      3891 => to_slv(opcode_type, 16#0E#),
      3892 => to_slv(opcode_type, 16#09#),
      3893 => to_slv(opcode_type, 16#08#),
      3894 => to_slv(opcode_type, 16#0B#),
      3895 => to_slv(opcode_type, 16#0C#),
      3896 => to_slv(opcode_type, 16#09#),
      3897 => to_slv(opcode_type, 16#0E#),
      3898 => to_slv(opcode_type, 16#0A#),
      3899 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#09#),
      3905 => to_slv(opcode_type, 16#09#),
      3906 => to_slv(opcode_type, 16#06#),
      3907 => to_slv(opcode_type, 16#08#),
      3908 => to_slv(opcode_type, 16#0F#),
      3909 => to_slv(opcode_type, 16#10#),
      3910 => to_slv(opcode_type, 16#08#),
      3911 => to_slv(opcode_type, 16#0E#),
      3912 => to_slv(opcode_type, 16#0D#),
      3913 => to_slv(opcode_type, 16#03#),
      3914 => to_slv(opcode_type, 16#05#),
      3915 => to_slv(opcode_type, 16#CE#),
      3916 => to_slv(opcode_type, 16#06#),
      3917 => to_slv(opcode_type, 16#07#),
      3918 => to_slv(opcode_type, 16#08#),
      3919 => to_slv(opcode_type, 16#0E#),
      3920 => to_slv(opcode_type, 16#61#),
      3921 => to_slv(opcode_type, 16#09#),
      3922 => to_slv(opcode_type, 16#0B#),
      3923 => to_slv(opcode_type, 16#11#),
      3924 => to_slv(opcode_type, 16#06#),
      3925 => to_slv(opcode_type, 16#09#),
      3926 => to_slv(opcode_type, 16#0E#),
      3927 => to_slv(opcode_type, 16#0F#),
      3928 => to_slv(opcode_type, 16#09#),
      3929 => to_slv(opcode_type, 16#11#),
      3930 => to_slv(opcode_type, 16#0F#),
      3931 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#07#),
      3937 => to_slv(opcode_type, 16#07#),
      3938 => to_slv(opcode_type, 16#04#),
      3939 => to_slv(opcode_type, 16#07#),
      3940 => to_slv(opcode_type, 16#0F#),
      3941 => to_slv(opcode_type, 16#10#),
      3942 => to_slv(opcode_type, 16#07#),
      3943 => to_slv(opcode_type, 16#01#),
      3944 => to_slv(opcode_type, 16#0E#),
      3945 => to_slv(opcode_type, 16#07#),
      3946 => to_slv(opcode_type, 16#0B#),
      3947 => to_slv(opcode_type, 16#38#),
      3948 => to_slv(opcode_type, 16#07#),
      3949 => to_slv(opcode_type, 16#06#),
      3950 => to_slv(opcode_type, 16#09#),
      3951 => to_slv(opcode_type, 16#0C#),
      3952 => to_slv(opcode_type, 16#0D#),
      3953 => to_slv(opcode_type, 16#06#),
      3954 => to_slv(opcode_type, 16#10#),
      3955 => to_slv(opcode_type, 16#11#),
      3956 => to_slv(opcode_type, 16#06#),
      3957 => to_slv(opcode_type, 16#07#),
      3958 => to_slv(opcode_type, 16#0D#),
      3959 => to_slv(opcode_type, 16#0E#),
      3960 => to_slv(opcode_type, 16#07#),
      3961 => to_slv(opcode_type, 16#0D#),
      3962 => to_slv(opcode_type, 16#10#),
      3963 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#08#),
      3969 => to_slv(opcode_type, 16#06#),
      3970 => to_slv(opcode_type, 16#08#),
      3971 => to_slv(opcode_type, 16#05#),
      3972 => to_slv(opcode_type, 16#0A#),
      3973 => to_slv(opcode_type, 16#02#),
      3974 => to_slv(opcode_type, 16#0D#),
      3975 => to_slv(opcode_type, 16#09#),
      3976 => to_slv(opcode_type, 16#06#),
      3977 => to_slv(opcode_type, 16#0E#),
      3978 => to_slv(opcode_type, 16#0A#),
      3979 => to_slv(opcode_type, 16#05#),
      3980 => to_slv(opcode_type, 16#11#),
      3981 => to_slv(opcode_type, 16#08#),
      3982 => to_slv(opcode_type, 16#08#),
      3983 => to_slv(opcode_type, 16#03#),
      3984 => to_slv(opcode_type, 16#0D#),
      3985 => to_slv(opcode_type, 16#09#),
      3986 => to_slv(opcode_type, 16#C3#),
      3987 => to_slv(opcode_type, 16#AF#),
      3988 => to_slv(opcode_type, 16#06#),
      3989 => to_slv(opcode_type, 16#08#),
      3990 => to_slv(opcode_type, 16#0D#),
      3991 => to_slv(opcode_type, 16#0F#),
      3992 => to_slv(opcode_type, 16#08#),
      3993 => to_slv(opcode_type, 16#0A#),
      3994 => to_slv(opcode_type, 16#11#),
      3995 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#07#),
      4001 => to_slv(opcode_type, 16#08#),
      4002 => to_slv(opcode_type, 16#02#),
      4003 => to_slv(opcode_type, 16#02#),
      4004 => to_slv(opcode_type, 16#0E#),
      4005 => to_slv(opcode_type, 16#06#),
      4006 => to_slv(opcode_type, 16#07#),
      4007 => to_slv(opcode_type, 16#0C#),
      4008 => to_slv(opcode_type, 16#11#),
      4009 => to_slv(opcode_type, 16#08#),
      4010 => to_slv(opcode_type, 16#10#),
      4011 => to_slv(opcode_type, 16#0D#),
      4012 => to_slv(opcode_type, 16#06#),
      4013 => to_slv(opcode_type, 16#08#),
      4014 => to_slv(opcode_type, 16#07#),
      4015 => to_slv(opcode_type, 16#0A#),
      4016 => to_slv(opcode_type, 16#0C#),
      4017 => to_slv(opcode_type, 16#08#),
      4018 => to_slv(opcode_type, 16#0B#),
      4019 => to_slv(opcode_type, 16#0B#),
      4020 => to_slv(opcode_type, 16#09#),
      4021 => to_slv(opcode_type, 16#08#),
      4022 => to_slv(opcode_type, 16#0A#),
      4023 => to_slv(opcode_type, 16#0F#),
      4024 => to_slv(opcode_type, 16#08#),
      4025 => to_slv(opcode_type, 16#0F#),
      4026 => to_slv(opcode_type, 16#0D#),
      4027 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#06#),
      4033 => to_slv(opcode_type, 16#06#),
      4034 => to_slv(opcode_type, 16#04#),
      4035 => to_slv(opcode_type, 16#07#),
      4036 => to_slv(opcode_type, 16#0B#),
      4037 => to_slv(opcode_type, 16#0E#),
      4038 => to_slv(opcode_type, 16#08#),
      4039 => to_slv(opcode_type, 16#08#),
      4040 => to_slv(opcode_type, 16#0D#),
      4041 => to_slv(opcode_type, 16#10#),
      4042 => to_slv(opcode_type, 16#08#),
      4043 => to_slv(opcode_type, 16#0D#),
      4044 => to_slv(opcode_type, 16#11#),
      4045 => to_slv(opcode_type, 16#09#),
      4046 => to_slv(opcode_type, 16#08#),
      4047 => to_slv(opcode_type, 16#05#),
      4048 => to_slv(opcode_type, 16#11#),
      4049 => to_slv(opcode_type, 16#07#),
      4050 => to_slv(opcode_type, 16#59#),
      4051 => to_slv(opcode_type, 16#0D#),
      4052 => to_slv(opcode_type, 16#06#),
      4053 => to_slv(opcode_type, 16#06#),
      4054 => to_slv(opcode_type, 16#0D#),
      4055 => to_slv(opcode_type, 16#10#),
      4056 => to_slv(opcode_type, 16#08#),
      4057 => to_slv(opcode_type, 16#0D#),
      4058 => to_slv(opcode_type, 16#0B#),
      4059 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#08#),
      4066 => to_slv(opcode_type, 16#04#),
      4067 => to_slv(opcode_type, 16#08#),
      4068 => to_slv(opcode_type, 16#0E#),
      4069 => to_slv(opcode_type, 16#0A#),
      4070 => to_slv(opcode_type, 16#07#),
      4071 => to_slv(opcode_type, 16#03#),
      4072 => to_slv(opcode_type, 16#96#),
      4073 => to_slv(opcode_type, 16#08#),
      4074 => to_slv(opcode_type, 16#0D#),
      4075 => to_slv(opcode_type, 16#0E#),
      4076 => to_slv(opcode_type, 16#09#),
      4077 => to_slv(opcode_type, 16#08#),
      4078 => to_slv(opcode_type, 16#06#),
      4079 => to_slv(opcode_type, 16#0C#),
      4080 => to_slv(opcode_type, 16#10#),
      4081 => to_slv(opcode_type, 16#07#),
      4082 => to_slv(opcode_type, 16#0C#),
      4083 => to_slv(opcode_type, 16#0C#),
      4084 => to_slv(opcode_type, 16#07#),
      4085 => to_slv(opcode_type, 16#08#),
      4086 => to_slv(opcode_type, 16#10#),
      4087 => to_slv(opcode_type, 16#0C#),
      4088 => to_slv(opcode_type, 16#09#),
      4089 => to_slv(opcode_type, 16#0A#),
      4090 => to_slv(opcode_type, 16#0B#),
      4091 to 4095 => (others => '0')
  ),

    -- Bin `28`...
    27 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#06#),
      1 => to_slv(opcode_type, 16#09#),
      2 => to_slv(opcode_type, 16#03#),
      3 => to_slv(opcode_type, 16#07#),
      4 => to_slv(opcode_type, 16#76#),
      5 => to_slv(opcode_type, 16#0D#),
      6 => to_slv(opcode_type, 16#06#),
      7 => to_slv(opcode_type, 16#09#),
      8 => to_slv(opcode_type, 16#0B#),
      9 => to_slv(opcode_type, 16#0C#),
      10 => to_slv(opcode_type, 16#07#),
      11 => to_slv(opcode_type, 16#B2#),
      12 => to_slv(opcode_type, 16#10#),
      13 => to_slv(opcode_type, 16#06#),
      14 => to_slv(opcode_type, 16#09#),
      15 => to_slv(opcode_type, 16#06#),
      16 => to_slv(opcode_type, 16#11#),
      17 => to_slv(opcode_type, 16#0C#),
      18 => to_slv(opcode_type, 16#06#),
      19 => to_slv(opcode_type, 16#0A#),
      20 => to_slv(opcode_type, 16#0A#),
      21 => to_slv(opcode_type, 16#06#),
      22 => to_slv(opcode_type, 16#06#),
      23 => to_slv(opcode_type, 16#0A#),
      24 => to_slv(opcode_type, 16#37#),
      25 => to_slv(opcode_type, 16#09#),
      26 => to_slv(opcode_type, 16#0C#),
      27 => to_slv(opcode_type, 16#11#),
      28 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#07#),
      33 => to_slv(opcode_type, 16#08#),
      34 => to_slv(opcode_type, 16#05#),
      35 => to_slv(opcode_type, 16#06#),
      36 => to_slv(opcode_type, 16#0A#),
      37 => to_slv(opcode_type, 16#0B#),
      38 => to_slv(opcode_type, 16#07#),
      39 => to_slv(opcode_type, 16#09#),
      40 => to_slv(opcode_type, 16#0B#),
      41 => to_slv(opcode_type, 16#0C#),
      42 => to_slv(opcode_type, 16#09#),
      43 => to_slv(opcode_type, 16#0C#),
      44 => to_slv(opcode_type, 16#0B#),
      45 => to_slv(opcode_type, 16#06#),
      46 => to_slv(opcode_type, 16#09#),
      47 => to_slv(opcode_type, 16#09#),
      48 => to_slv(opcode_type, 16#0D#),
      49 => to_slv(opcode_type, 16#10#),
      50 => to_slv(opcode_type, 16#08#),
      51 => to_slv(opcode_type, 16#0B#),
      52 => to_slv(opcode_type, 16#0D#),
      53 => to_slv(opcode_type, 16#09#),
      54 => to_slv(opcode_type, 16#08#),
      55 => to_slv(opcode_type, 16#E7#),
      56 => to_slv(opcode_type, 16#0A#),
      57 => to_slv(opcode_type, 16#08#),
      58 => to_slv(opcode_type, 16#0A#),
      59 => to_slv(opcode_type, 16#0B#),
      60 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#09#),
      65 => to_slv(opcode_type, 16#08#),
      66 => to_slv(opcode_type, 16#05#),
      67 => to_slv(opcode_type, 16#08#),
      68 => to_slv(opcode_type, 16#0E#),
      69 => to_slv(opcode_type, 16#0B#),
      70 => to_slv(opcode_type, 16#06#),
      71 => to_slv(opcode_type, 16#09#),
      72 => to_slv(opcode_type, 16#11#),
      73 => to_slv(opcode_type, 16#C7#),
      74 => to_slv(opcode_type, 16#08#),
      75 => to_slv(opcode_type, 16#0C#),
      76 => to_slv(opcode_type, 16#0F#),
      77 => to_slv(opcode_type, 16#08#),
      78 => to_slv(opcode_type, 16#06#),
      79 => to_slv(opcode_type, 16#07#),
      80 => to_slv(opcode_type, 16#11#),
      81 => to_slv(opcode_type, 16#0A#),
      82 => to_slv(opcode_type, 16#07#),
      83 => to_slv(opcode_type, 16#0C#),
      84 => to_slv(opcode_type, 16#11#),
      85 => to_slv(opcode_type, 16#06#),
      86 => to_slv(opcode_type, 16#07#),
      87 => to_slv(opcode_type, 16#0A#),
      88 => to_slv(opcode_type, 16#0B#),
      89 => to_slv(opcode_type, 16#06#),
      90 => to_slv(opcode_type, 16#0B#),
      91 => to_slv(opcode_type, 16#11#),
      92 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#08#),
      97 => to_slv(opcode_type, 16#07#),
      98 => to_slv(opcode_type, 16#01#),
      99 => to_slv(opcode_type, 16#08#),
      100 => to_slv(opcode_type, 16#10#),
      101 => to_slv(opcode_type, 16#0B#),
      102 => to_slv(opcode_type, 16#08#),
      103 => to_slv(opcode_type, 16#07#),
      104 => to_slv(opcode_type, 16#0B#),
      105 => to_slv(opcode_type, 16#0A#),
      106 => to_slv(opcode_type, 16#08#),
      107 => to_slv(opcode_type, 16#0D#),
      108 => to_slv(opcode_type, 16#0F#),
      109 => to_slv(opcode_type, 16#07#),
      110 => to_slv(opcode_type, 16#07#),
      111 => to_slv(opcode_type, 16#06#),
      112 => to_slv(opcode_type, 16#0D#),
      113 => to_slv(opcode_type, 16#11#),
      114 => to_slv(opcode_type, 16#08#),
      115 => to_slv(opcode_type, 16#0C#),
      116 => to_slv(opcode_type, 16#0E#),
      117 => to_slv(opcode_type, 16#08#),
      118 => to_slv(opcode_type, 16#06#),
      119 => to_slv(opcode_type, 16#9A#),
      120 => to_slv(opcode_type, 16#0B#),
      121 => to_slv(opcode_type, 16#06#),
      122 => to_slv(opcode_type, 16#0E#),
      123 => to_slv(opcode_type, 16#0D#),
      124 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#08#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#07#),
      131 => to_slv(opcode_type, 16#03#),
      132 => to_slv(opcode_type, 16#11#),
      133 => to_slv(opcode_type, 16#03#),
      134 => to_slv(opcode_type, 16#11#),
      135 => to_slv(opcode_type, 16#08#),
      136 => to_slv(opcode_type, 16#05#),
      137 => to_slv(opcode_type, 16#43#),
      138 => to_slv(opcode_type, 16#08#),
      139 => to_slv(opcode_type, 16#0D#),
      140 => to_slv(opcode_type, 16#0B#),
      141 => to_slv(opcode_type, 16#09#),
      142 => to_slv(opcode_type, 16#08#),
      143 => to_slv(opcode_type, 16#06#),
      144 => to_slv(opcode_type, 16#38#),
      145 => to_slv(opcode_type, 16#0F#),
      146 => to_slv(opcode_type, 16#09#),
      147 => to_slv(opcode_type, 16#0F#),
      148 => to_slv(opcode_type, 16#0F#),
      149 => to_slv(opcode_type, 16#06#),
      150 => to_slv(opcode_type, 16#09#),
      151 => to_slv(opcode_type, 16#0C#),
      152 => to_slv(opcode_type, 16#0F#),
      153 => to_slv(opcode_type, 16#08#),
      154 => to_slv(opcode_type, 16#0C#),
      155 => to_slv(opcode_type, 16#11#),
      156 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#07#),
      161 => to_slv(opcode_type, 16#06#),
      162 => to_slv(opcode_type, 16#07#),
      163 => to_slv(opcode_type, 16#09#),
      164 => to_slv(opcode_type, 16#0C#),
      165 => to_slv(opcode_type, 16#0E#),
      166 => to_slv(opcode_type, 16#08#),
      167 => to_slv(opcode_type, 16#0B#),
      168 => to_slv(opcode_type, 16#0B#),
      169 => to_slv(opcode_type, 16#02#),
      170 => to_slv(opcode_type, 16#08#),
      171 => to_slv(opcode_type, 16#0F#),
      172 => to_slv(opcode_type, 16#0C#),
      173 => to_slv(opcode_type, 16#09#),
      174 => to_slv(opcode_type, 16#08#),
      175 => to_slv(opcode_type, 16#09#),
      176 => to_slv(opcode_type, 16#0B#),
      177 => to_slv(opcode_type, 16#0F#),
      178 => to_slv(opcode_type, 16#06#),
      179 => to_slv(opcode_type, 16#0B#),
      180 => to_slv(opcode_type, 16#0D#),
      181 => to_slv(opcode_type, 16#09#),
      182 => to_slv(opcode_type, 16#08#),
      183 => to_slv(opcode_type, 16#0E#),
      184 => to_slv(opcode_type, 16#0D#),
      185 => to_slv(opcode_type, 16#07#),
      186 => to_slv(opcode_type, 16#0E#),
      187 => to_slv(opcode_type, 16#0B#),
      188 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#06#),
      193 => to_slv(opcode_type, 16#06#),
      194 => to_slv(opcode_type, 16#08#),
      195 => to_slv(opcode_type, 16#05#),
      196 => to_slv(opcode_type, 16#3C#),
      197 => to_slv(opcode_type, 16#09#),
      198 => to_slv(opcode_type, 16#10#),
      199 => to_slv(opcode_type, 16#0E#),
      200 => to_slv(opcode_type, 16#08#),
      201 => to_slv(opcode_type, 16#02#),
      202 => to_slv(opcode_type, 16#11#),
      203 => to_slv(opcode_type, 16#01#),
      204 => to_slv(opcode_type, 16#0D#),
      205 => to_slv(opcode_type, 16#08#),
      206 => to_slv(opcode_type, 16#06#),
      207 => to_slv(opcode_type, 16#07#),
      208 => to_slv(opcode_type, 16#55#),
      209 => to_slv(opcode_type, 16#11#),
      210 => to_slv(opcode_type, 16#08#),
      211 => to_slv(opcode_type, 16#C7#),
      212 => to_slv(opcode_type, 16#0F#),
      213 => to_slv(opcode_type, 16#09#),
      214 => to_slv(opcode_type, 16#08#),
      215 => to_slv(opcode_type, 16#11#),
      216 => to_slv(opcode_type, 16#0B#),
      217 => to_slv(opcode_type, 16#06#),
      218 => to_slv(opcode_type, 16#0C#),
      219 => to_slv(opcode_type, 16#0F#),
      220 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#08#),
      225 => to_slv(opcode_type, 16#06#),
      226 => to_slv(opcode_type, 16#09#),
      227 => to_slv(opcode_type, 16#03#),
      228 => to_slv(opcode_type, 16#0A#),
      229 => to_slv(opcode_type, 16#07#),
      230 => to_slv(opcode_type, 16#11#),
      231 => to_slv(opcode_type, 16#0F#),
      232 => to_slv(opcode_type, 16#07#),
      233 => to_slv(opcode_type, 16#01#),
      234 => to_slv(opcode_type, 16#0F#),
      235 => to_slv(opcode_type, 16#07#),
      236 => to_slv(opcode_type, 16#0C#),
      237 => to_slv(opcode_type, 16#0D#),
      238 => to_slv(opcode_type, 16#06#),
      239 => to_slv(opcode_type, 16#06#),
      240 => to_slv(opcode_type, 16#04#),
      241 => to_slv(opcode_type, 16#0B#),
      242 => to_slv(opcode_type, 16#09#),
      243 => to_slv(opcode_type, 16#0A#),
      244 => to_slv(opcode_type, 16#0F#),
      245 => to_slv(opcode_type, 16#06#),
      246 => to_slv(opcode_type, 16#07#),
      247 => to_slv(opcode_type, 16#0B#),
      248 => to_slv(opcode_type, 16#0B#),
      249 => to_slv(opcode_type, 16#09#),
      250 => to_slv(opcode_type, 16#0E#),
      251 => to_slv(opcode_type, 16#0A#),
      252 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#06#),
      257 => to_slv(opcode_type, 16#08#),
      258 => to_slv(opcode_type, 16#06#),
      259 => to_slv(opcode_type, 16#06#),
      260 => to_slv(opcode_type, 16#0C#),
      261 => to_slv(opcode_type, 16#0D#),
      262 => to_slv(opcode_type, 16#02#),
      263 => to_slv(opcode_type, 16#0E#),
      264 => to_slv(opcode_type, 16#09#),
      265 => to_slv(opcode_type, 16#06#),
      266 => to_slv(opcode_type, 16#0D#),
      267 => to_slv(opcode_type, 16#0E#),
      268 => to_slv(opcode_type, 16#03#),
      269 => to_slv(opcode_type, 16#11#),
      270 => to_slv(opcode_type, 16#07#),
      271 => to_slv(opcode_type, 16#07#),
      272 => to_slv(opcode_type, 16#09#),
      273 => to_slv(opcode_type, 16#0D#),
      274 => to_slv(opcode_type, 16#11#),
      275 => to_slv(opcode_type, 16#01#),
      276 => to_slv(opcode_type, 16#11#),
      277 => to_slv(opcode_type, 16#07#),
      278 => to_slv(opcode_type, 16#08#),
      279 => to_slv(opcode_type, 16#10#),
      280 => to_slv(opcode_type, 16#10#),
      281 => to_slv(opcode_type, 16#09#),
      282 => to_slv(opcode_type, 16#0A#),
      283 => to_slv(opcode_type, 16#0F#),
      284 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#09#),
      289 => to_slv(opcode_type, 16#07#),
      290 => to_slv(opcode_type, 16#08#),
      291 => to_slv(opcode_type, 16#06#),
      292 => to_slv(opcode_type, 16#0C#),
      293 => to_slv(opcode_type, 16#0D#),
      294 => to_slv(opcode_type, 16#07#),
      295 => to_slv(opcode_type, 16#0C#),
      296 => to_slv(opcode_type, 16#0A#),
      297 => to_slv(opcode_type, 16#06#),
      298 => to_slv(opcode_type, 16#02#),
      299 => to_slv(opcode_type, 16#0A#),
      300 => to_slv(opcode_type, 16#03#),
      301 => to_slv(opcode_type, 16#11#),
      302 => to_slv(opcode_type, 16#09#),
      303 => to_slv(opcode_type, 16#07#),
      304 => to_slv(opcode_type, 16#07#),
      305 => to_slv(opcode_type, 16#A5#),
      306 => to_slv(opcode_type, 16#0A#),
      307 => to_slv(opcode_type, 16#09#),
      308 => to_slv(opcode_type, 16#10#),
      309 => to_slv(opcode_type, 16#11#),
      310 => to_slv(opcode_type, 16#09#),
      311 => to_slv(opcode_type, 16#04#),
      312 => to_slv(opcode_type, 16#10#),
      313 => to_slv(opcode_type, 16#07#),
      314 => to_slv(opcode_type, 16#36#),
      315 => to_slv(opcode_type, 16#0B#),
      316 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#06#),
      321 => to_slv(opcode_type, 16#07#),
      322 => to_slv(opcode_type, 16#04#),
      323 => to_slv(opcode_type, 16#06#),
      324 => to_slv(opcode_type, 16#0F#),
      325 => to_slv(opcode_type, 16#0A#),
      326 => to_slv(opcode_type, 16#07#),
      327 => to_slv(opcode_type, 16#08#),
      328 => to_slv(opcode_type, 16#88#),
      329 => to_slv(opcode_type, 16#0A#),
      330 => to_slv(opcode_type, 16#07#),
      331 => to_slv(opcode_type, 16#0B#),
      332 => to_slv(opcode_type, 16#0A#),
      333 => to_slv(opcode_type, 16#08#),
      334 => to_slv(opcode_type, 16#07#),
      335 => to_slv(opcode_type, 16#08#),
      336 => to_slv(opcode_type, 16#0C#),
      337 => to_slv(opcode_type, 16#0A#),
      338 => to_slv(opcode_type, 16#08#),
      339 => to_slv(opcode_type, 16#15#),
      340 => to_slv(opcode_type, 16#0B#),
      341 => to_slv(opcode_type, 16#08#),
      342 => to_slv(opcode_type, 16#06#),
      343 => to_slv(opcode_type, 16#11#),
      344 => to_slv(opcode_type, 16#0F#),
      345 => to_slv(opcode_type, 16#08#),
      346 => to_slv(opcode_type, 16#BF#),
      347 => to_slv(opcode_type, 16#0E#),
      348 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#07#),
      353 => to_slv(opcode_type, 16#06#),
      354 => to_slv(opcode_type, 16#02#),
      355 => to_slv(opcode_type, 16#06#),
      356 => to_slv(opcode_type, 16#0A#),
      357 => to_slv(opcode_type, 16#10#),
      358 => to_slv(opcode_type, 16#08#),
      359 => to_slv(opcode_type, 16#08#),
      360 => to_slv(opcode_type, 16#0A#),
      361 => to_slv(opcode_type, 16#0D#),
      362 => to_slv(opcode_type, 16#06#),
      363 => to_slv(opcode_type, 16#0E#),
      364 => to_slv(opcode_type, 16#0D#),
      365 => to_slv(opcode_type, 16#09#),
      366 => to_slv(opcode_type, 16#06#),
      367 => to_slv(opcode_type, 16#06#),
      368 => to_slv(opcode_type, 16#0D#),
      369 => to_slv(opcode_type, 16#0F#),
      370 => to_slv(opcode_type, 16#08#),
      371 => to_slv(opcode_type, 16#0A#),
      372 => to_slv(opcode_type, 16#0B#),
      373 => to_slv(opcode_type, 16#07#),
      374 => to_slv(opcode_type, 16#07#),
      375 => to_slv(opcode_type, 16#0F#),
      376 => to_slv(opcode_type, 16#0A#),
      377 => to_slv(opcode_type, 16#07#),
      378 => to_slv(opcode_type, 16#0C#),
      379 => to_slv(opcode_type, 16#0F#),
      380 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#08#),
      385 => to_slv(opcode_type, 16#06#),
      386 => to_slv(opcode_type, 16#05#),
      387 => to_slv(opcode_type, 16#09#),
      388 => to_slv(opcode_type, 16#10#),
      389 => to_slv(opcode_type, 16#30#),
      390 => to_slv(opcode_type, 16#07#),
      391 => to_slv(opcode_type, 16#07#),
      392 => to_slv(opcode_type, 16#EE#),
      393 => to_slv(opcode_type, 16#11#),
      394 => to_slv(opcode_type, 16#08#),
      395 => to_slv(opcode_type, 16#10#),
      396 => to_slv(opcode_type, 16#A1#),
      397 => to_slv(opcode_type, 16#07#),
      398 => to_slv(opcode_type, 16#06#),
      399 => to_slv(opcode_type, 16#08#),
      400 => to_slv(opcode_type, 16#0B#),
      401 => to_slv(opcode_type, 16#0F#),
      402 => to_slv(opcode_type, 16#06#),
      403 => to_slv(opcode_type, 16#10#),
      404 => to_slv(opcode_type, 16#0F#),
      405 => to_slv(opcode_type, 16#06#),
      406 => to_slv(opcode_type, 16#08#),
      407 => to_slv(opcode_type, 16#0D#),
      408 => to_slv(opcode_type, 16#10#),
      409 => to_slv(opcode_type, 16#08#),
      410 => to_slv(opcode_type, 16#0C#),
      411 => to_slv(opcode_type, 16#11#),
      412 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#06#),
      417 => to_slv(opcode_type, 16#09#),
      418 => to_slv(opcode_type, 16#09#),
      419 => to_slv(opcode_type, 16#07#),
      420 => to_slv(opcode_type, 16#0C#),
      421 => to_slv(opcode_type, 16#0A#),
      422 => to_slv(opcode_type, 16#05#),
      423 => to_slv(opcode_type, 16#D3#),
      424 => to_slv(opcode_type, 16#07#),
      425 => to_slv(opcode_type, 16#03#),
      426 => to_slv(opcode_type, 16#10#),
      427 => to_slv(opcode_type, 16#09#),
      428 => to_slv(opcode_type, 16#10#),
      429 => to_slv(opcode_type, 16#C0#),
      430 => to_slv(opcode_type, 16#08#),
      431 => to_slv(opcode_type, 16#09#),
      432 => to_slv(opcode_type, 16#07#),
      433 => to_slv(opcode_type, 16#4A#),
      434 => to_slv(opcode_type, 16#11#),
      435 => to_slv(opcode_type, 16#01#),
      436 => to_slv(opcode_type, 16#10#),
      437 => to_slv(opcode_type, 16#09#),
      438 => to_slv(opcode_type, 16#09#),
      439 => to_slv(opcode_type, 16#0D#),
      440 => to_slv(opcode_type, 16#0F#),
      441 => to_slv(opcode_type, 16#08#),
      442 => to_slv(opcode_type, 16#7D#),
      443 => to_slv(opcode_type, 16#0F#),
      444 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#09#),
      449 => to_slv(opcode_type, 16#09#),
      450 => to_slv(opcode_type, 16#09#),
      451 => to_slv(opcode_type, 16#01#),
      452 => to_slv(opcode_type, 16#0A#),
      453 => to_slv(opcode_type, 16#03#),
      454 => to_slv(opcode_type, 16#0E#),
      455 => to_slv(opcode_type, 16#09#),
      456 => to_slv(opcode_type, 16#08#),
      457 => to_slv(opcode_type, 16#10#),
      458 => to_slv(opcode_type, 16#0D#),
      459 => to_slv(opcode_type, 16#07#),
      460 => to_slv(opcode_type, 16#0B#),
      461 => to_slv(opcode_type, 16#45#),
      462 => to_slv(opcode_type, 16#09#),
      463 => to_slv(opcode_type, 16#09#),
      464 => to_slv(opcode_type, 16#04#),
      465 => to_slv(opcode_type, 16#11#),
      466 => to_slv(opcode_type, 16#08#),
      467 => to_slv(opcode_type, 16#11#),
      468 => to_slv(opcode_type, 16#0F#),
      469 => to_slv(opcode_type, 16#06#),
      470 => to_slv(opcode_type, 16#06#),
      471 => to_slv(opcode_type, 16#0E#),
      472 => to_slv(opcode_type, 16#11#),
      473 => to_slv(opcode_type, 16#06#),
      474 => to_slv(opcode_type, 16#0B#),
      475 => to_slv(opcode_type, 16#0D#),
      476 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#07#),
      481 => to_slv(opcode_type, 16#08#),
      482 => to_slv(opcode_type, 16#08#),
      483 => to_slv(opcode_type, 16#03#),
      484 => to_slv(opcode_type, 16#0B#),
      485 => to_slv(opcode_type, 16#01#),
      486 => to_slv(opcode_type, 16#E1#),
      487 => to_slv(opcode_type, 16#07#),
      488 => to_slv(opcode_type, 16#04#),
      489 => to_slv(opcode_type, 16#0D#),
      490 => to_slv(opcode_type, 16#06#),
      491 => to_slv(opcode_type, 16#0A#),
      492 => to_slv(opcode_type, 16#0D#),
      493 => to_slv(opcode_type, 16#06#),
      494 => to_slv(opcode_type, 16#07#),
      495 => to_slv(opcode_type, 16#08#),
      496 => to_slv(opcode_type, 16#11#),
      497 => to_slv(opcode_type, 16#11#),
      498 => to_slv(opcode_type, 16#09#),
      499 => to_slv(opcode_type, 16#0F#),
      500 => to_slv(opcode_type, 16#0D#),
      501 => to_slv(opcode_type, 16#07#),
      502 => to_slv(opcode_type, 16#09#),
      503 => to_slv(opcode_type, 16#0B#),
      504 => to_slv(opcode_type, 16#11#),
      505 => to_slv(opcode_type, 16#07#),
      506 => to_slv(opcode_type, 16#CB#),
      507 => to_slv(opcode_type, 16#10#),
      508 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#07#),
      513 => to_slv(opcode_type, 16#06#),
      514 => to_slv(opcode_type, 16#06#),
      515 => to_slv(opcode_type, 16#02#),
      516 => to_slv(opcode_type, 16#11#),
      517 => to_slv(opcode_type, 16#08#),
      518 => to_slv(opcode_type, 16#0A#),
      519 => to_slv(opcode_type, 16#0E#),
      520 => to_slv(opcode_type, 16#09#),
      521 => to_slv(opcode_type, 16#09#),
      522 => to_slv(opcode_type, 16#A5#),
      523 => to_slv(opcode_type, 16#0C#),
      524 => to_slv(opcode_type, 16#03#),
      525 => to_slv(opcode_type, 16#11#),
      526 => to_slv(opcode_type, 16#07#),
      527 => to_slv(opcode_type, 16#07#),
      528 => to_slv(opcode_type, 16#05#),
      529 => to_slv(opcode_type, 16#9A#),
      530 => to_slv(opcode_type, 16#07#),
      531 => to_slv(opcode_type, 16#0D#),
      532 => to_slv(opcode_type, 16#0B#),
      533 => to_slv(opcode_type, 16#09#),
      534 => to_slv(opcode_type, 16#06#),
      535 => to_slv(opcode_type, 16#2F#),
      536 => to_slv(opcode_type, 16#10#),
      537 => to_slv(opcode_type, 16#07#),
      538 => to_slv(opcode_type, 16#92#),
      539 => to_slv(opcode_type, 16#0C#),
      540 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#08#),
      545 => to_slv(opcode_type, 16#07#),
      546 => to_slv(opcode_type, 16#09#),
      547 => to_slv(opcode_type, 16#03#),
      548 => to_slv(opcode_type, 16#0F#),
      549 => to_slv(opcode_type, 16#01#),
      550 => to_slv(opcode_type, 16#0B#),
      551 => to_slv(opcode_type, 16#07#),
      552 => to_slv(opcode_type, 16#08#),
      553 => to_slv(opcode_type, 16#0B#),
      554 => to_slv(opcode_type, 16#0F#),
      555 => to_slv(opcode_type, 16#01#),
      556 => to_slv(opcode_type, 16#0F#),
      557 => to_slv(opcode_type, 16#08#),
      558 => to_slv(opcode_type, 16#09#),
      559 => to_slv(opcode_type, 16#07#),
      560 => to_slv(opcode_type, 16#0F#),
      561 => to_slv(opcode_type, 16#32#),
      562 => to_slv(opcode_type, 16#07#),
      563 => to_slv(opcode_type, 16#0E#),
      564 => to_slv(opcode_type, 16#0E#),
      565 => to_slv(opcode_type, 16#08#),
      566 => to_slv(opcode_type, 16#09#),
      567 => to_slv(opcode_type, 16#50#),
      568 => to_slv(opcode_type, 16#11#),
      569 => to_slv(opcode_type, 16#09#),
      570 => to_slv(opcode_type, 16#0B#),
      571 => to_slv(opcode_type, 16#10#),
      572 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#07#),
      577 => to_slv(opcode_type, 16#07#),
      578 => to_slv(opcode_type, 16#09#),
      579 => to_slv(opcode_type, 16#04#),
      580 => to_slv(opcode_type, 16#0A#),
      581 => to_slv(opcode_type, 16#09#),
      582 => to_slv(opcode_type, 16#0A#),
      583 => to_slv(opcode_type, 16#0E#),
      584 => to_slv(opcode_type, 16#09#),
      585 => to_slv(opcode_type, 16#01#),
      586 => to_slv(opcode_type, 16#10#),
      587 => to_slv(opcode_type, 16#07#),
      588 => to_slv(opcode_type, 16#11#),
      589 => to_slv(opcode_type, 16#10#),
      590 => to_slv(opcode_type, 16#09#),
      591 => to_slv(opcode_type, 16#06#),
      592 => to_slv(opcode_type, 16#09#),
      593 => to_slv(opcode_type, 16#10#),
      594 => to_slv(opcode_type, 16#0F#),
      595 => to_slv(opcode_type, 16#03#),
      596 => to_slv(opcode_type, 16#11#),
      597 => to_slv(opcode_type, 16#07#),
      598 => to_slv(opcode_type, 16#07#),
      599 => to_slv(opcode_type, 16#0A#),
      600 => to_slv(opcode_type, 16#0C#),
      601 => to_slv(opcode_type, 16#07#),
      602 => to_slv(opcode_type, 16#E3#),
      603 => to_slv(opcode_type, 16#0A#),
      604 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#09#),
      609 => to_slv(opcode_type, 16#09#),
      610 => to_slv(opcode_type, 16#05#),
      611 => to_slv(opcode_type, 16#08#),
      612 => to_slv(opcode_type, 16#0B#),
      613 => to_slv(opcode_type, 16#10#),
      614 => to_slv(opcode_type, 16#08#),
      615 => to_slv(opcode_type, 16#08#),
      616 => to_slv(opcode_type, 16#0B#),
      617 => to_slv(opcode_type, 16#0A#),
      618 => to_slv(opcode_type, 16#08#),
      619 => to_slv(opcode_type, 16#0E#),
      620 => to_slv(opcode_type, 16#10#),
      621 => to_slv(opcode_type, 16#09#),
      622 => to_slv(opcode_type, 16#06#),
      623 => to_slv(opcode_type, 16#09#),
      624 => to_slv(opcode_type, 16#3B#),
      625 => to_slv(opcode_type, 16#11#),
      626 => to_slv(opcode_type, 16#07#),
      627 => to_slv(opcode_type, 16#10#),
      628 => to_slv(opcode_type, 16#10#),
      629 => to_slv(opcode_type, 16#08#),
      630 => to_slv(opcode_type, 16#06#),
      631 => to_slv(opcode_type, 16#0B#),
      632 => to_slv(opcode_type, 16#0E#),
      633 => to_slv(opcode_type, 16#07#),
      634 => to_slv(opcode_type, 16#0A#),
      635 => to_slv(opcode_type, 16#0A#),
      636 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#06#),
      641 => to_slv(opcode_type, 16#09#),
      642 => to_slv(opcode_type, 16#08#),
      643 => to_slv(opcode_type, 16#06#),
      644 => to_slv(opcode_type, 16#0E#),
      645 => to_slv(opcode_type, 16#0B#),
      646 => to_slv(opcode_type, 16#02#),
      647 => to_slv(opcode_type, 16#10#),
      648 => to_slv(opcode_type, 16#07#),
      649 => to_slv(opcode_type, 16#01#),
      650 => to_slv(opcode_type, 16#0F#),
      651 => to_slv(opcode_type, 16#08#),
      652 => to_slv(opcode_type, 16#10#),
      653 => to_slv(opcode_type, 16#0A#),
      654 => to_slv(opcode_type, 16#08#),
      655 => to_slv(opcode_type, 16#08#),
      656 => to_slv(opcode_type, 16#06#),
      657 => to_slv(opcode_type, 16#0C#),
      658 => to_slv(opcode_type, 16#0C#),
      659 => to_slv(opcode_type, 16#05#),
      660 => to_slv(opcode_type, 16#11#),
      661 => to_slv(opcode_type, 16#06#),
      662 => to_slv(opcode_type, 16#09#),
      663 => to_slv(opcode_type, 16#0C#),
      664 => to_slv(opcode_type, 16#0E#),
      665 => to_slv(opcode_type, 16#09#),
      666 => to_slv(opcode_type, 16#0B#),
      667 => to_slv(opcode_type, 16#0B#),
      668 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#09#),
      673 => to_slv(opcode_type, 16#08#),
      674 => to_slv(opcode_type, 16#06#),
      675 => to_slv(opcode_type, 16#01#),
      676 => to_slv(opcode_type, 16#0C#),
      677 => to_slv(opcode_type, 16#06#),
      678 => to_slv(opcode_type, 16#0F#),
      679 => to_slv(opcode_type, 16#0A#),
      680 => to_slv(opcode_type, 16#06#),
      681 => to_slv(opcode_type, 16#03#),
      682 => to_slv(opcode_type, 16#0E#),
      683 => to_slv(opcode_type, 16#07#),
      684 => to_slv(opcode_type, 16#0B#),
      685 => to_slv(opcode_type, 16#0C#),
      686 => to_slv(opcode_type, 16#06#),
      687 => to_slv(opcode_type, 16#06#),
      688 => to_slv(opcode_type, 16#07#),
      689 => to_slv(opcode_type, 16#0B#),
      690 => to_slv(opcode_type, 16#0C#),
      691 => to_slv(opcode_type, 16#01#),
      692 => to_slv(opcode_type, 16#0C#),
      693 => to_slv(opcode_type, 16#06#),
      694 => to_slv(opcode_type, 16#07#),
      695 => to_slv(opcode_type, 16#0A#),
      696 => to_slv(opcode_type, 16#11#),
      697 => to_slv(opcode_type, 16#07#),
      698 => to_slv(opcode_type, 16#0E#),
      699 => to_slv(opcode_type, 16#0F#),
      700 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#06#),
      705 => to_slv(opcode_type, 16#07#),
      706 => to_slv(opcode_type, 16#05#),
      707 => to_slv(opcode_type, 16#08#),
      708 => to_slv(opcode_type, 16#0E#),
      709 => to_slv(opcode_type, 16#0C#),
      710 => to_slv(opcode_type, 16#09#),
      711 => to_slv(opcode_type, 16#08#),
      712 => to_slv(opcode_type, 16#0F#),
      713 => to_slv(opcode_type, 16#10#),
      714 => to_slv(opcode_type, 16#08#),
      715 => to_slv(opcode_type, 16#10#),
      716 => to_slv(opcode_type, 16#0F#),
      717 => to_slv(opcode_type, 16#08#),
      718 => to_slv(opcode_type, 16#08#),
      719 => to_slv(opcode_type, 16#07#),
      720 => to_slv(opcode_type, 16#B9#),
      721 => to_slv(opcode_type, 16#0B#),
      722 => to_slv(opcode_type, 16#06#),
      723 => to_slv(opcode_type, 16#0D#),
      724 => to_slv(opcode_type, 16#10#),
      725 => to_slv(opcode_type, 16#07#),
      726 => to_slv(opcode_type, 16#06#),
      727 => to_slv(opcode_type, 16#0F#),
      728 => to_slv(opcode_type, 16#0F#),
      729 => to_slv(opcode_type, 16#08#),
      730 => to_slv(opcode_type, 16#0E#),
      731 => to_slv(opcode_type, 16#0A#),
      732 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#08#),
      737 => to_slv(opcode_type, 16#08#),
      738 => to_slv(opcode_type, 16#05#),
      739 => to_slv(opcode_type, 16#07#),
      740 => to_slv(opcode_type, 16#6B#),
      741 => to_slv(opcode_type, 16#CC#),
      742 => to_slv(opcode_type, 16#07#),
      743 => to_slv(opcode_type, 16#06#),
      744 => to_slv(opcode_type, 16#0B#),
      745 => to_slv(opcode_type, 16#11#),
      746 => to_slv(opcode_type, 16#08#),
      747 => to_slv(opcode_type, 16#0F#),
      748 => to_slv(opcode_type, 16#10#),
      749 => to_slv(opcode_type, 16#07#),
      750 => to_slv(opcode_type, 16#09#),
      751 => to_slv(opcode_type, 16#09#),
      752 => to_slv(opcode_type, 16#0F#),
      753 => to_slv(opcode_type, 16#0C#),
      754 => to_slv(opcode_type, 16#07#),
      755 => to_slv(opcode_type, 16#0E#),
      756 => to_slv(opcode_type, 16#E4#),
      757 => to_slv(opcode_type, 16#09#),
      758 => to_slv(opcode_type, 16#07#),
      759 => to_slv(opcode_type, 16#0A#),
      760 => to_slv(opcode_type, 16#0F#),
      761 => to_slv(opcode_type, 16#09#),
      762 => to_slv(opcode_type, 16#0E#),
      763 => to_slv(opcode_type, 16#10#),
      764 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#07#),
      769 => to_slv(opcode_type, 16#07#),
      770 => to_slv(opcode_type, 16#07#),
      771 => to_slv(opcode_type, 16#09#),
      772 => to_slv(opcode_type, 16#11#),
      773 => to_slv(opcode_type, 16#0E#),
      774 => to_slv(opcode_type, 16#05#),
      775 => to_slv(opcode_type, 16#0F#),
      776 => to_slv(opcode_type, 16#07#),
      777 => to_slv(opcode_type, 16#06#),
      778 => to_slv(opcode_type, 16#0B#),
      779 => to_slv(opcode_type, 16#10#),
      780 => to_slv(opcode_type, 16#06#),
      781 => to_slv(opcode_type, 16#11#),
      782 => to_slv(opcode_type, 16#10#),
      783 => to_slv(opcode_type, 16#09#),
      784 => to_slv(opcode_type, 16#06#),
      785 => to_slv(opcode_type, 16#07#),
      786 => to_slv(opcode_type, 16#0D#),
      787 => to_slv(opcode_type, 16#0D#),
      788 => to_slv(opcode_type, 16#01#),
      789 => to_slv(opcode_type, 16#11#),
      790 => to_slv(opcode_type, 16#09#),
      791 => to_slv(opcode_type, 16#06#),
      792 => to_slv(opcode_type, 16#0E#),
      793 => to_slv(opcode_type, 16#0C#),
      794 => to_slv(opcode_type, 16#02#),
      795 => to_slv(opcode_type, 16#0F#),
      796 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#07#),
      801 => to_slv(opcode_type, 16#09#),
      802 => to_slv(opcode_type, 16#01#),
      803 => to_slv(opcode_type, 16#09#),
      804 => to_slv(opcode_type, 16#0B#),
      805 => to_slv(opcode_type, 16#0B#),
      806 => to_slv(opcode_type, 16#09#),
      807 => to_slv(opcode_type, 16#07#),
      808 => to_slv(opcode_type, 16#0F#),
      809 => to_slv(opcode_type, 16#0F#),
      810 => to_slv(opcode_type, 16#06#),
      811 => to_slv(opcode_type, 16#0C#),
      812 => to_slv(opcode_type, 16#0C#),
      813 => to_slv(opcode_type, 16#07#),
      814 => to_slv(opcode_type, 16#06#),
      815 => to_slv(opcode_type, 16#07#),
      816 => to_slv(opcode_type, 16#0A#),
      817 => to_slv(opcode_type, 16#0C#),
      818 => to_slv(opcode_type, 16#07#),
      819 => to_slv(opcode_type, 16#11#),
      820 => to_slv(opcode_type, 16#0F#),
      821 => to_slv(opcode_type, 16#08#),
      822 => to_slv(opcode_type, 16#08#),
      823 => to_slv(opcode_type, 16#F6#),
      824 => to_slv(opcode_type, 16#0C#),
      825 => to_slv(opcode_type, 16#09#),
      826 => to_slv(opcode_type, 16#0F#),
      827 => to_slv(opcode_type, 16#8A#),
      828 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#06#),
      833 => to_slv(opcode_type, 16#06#),
      834 => to_slv(opcode_type, 16#05#),
      835 => to_slv(opcode_type, 16#07#),
      836 => to_slv(opcode_type, 16#0C#),
      837 => to_slv(opcode_type, 16#0D#),
      838 => to_slv(opcode_type, 16#09#),
      839 => to_slv(opcode_type, 16#07#),
      840 => to_slv(opcode_type, 16#10#),
      841 => to_slv(opcode_type, 16#0F#),
      842 => to_slv(opcode_type, 16#09#),
      843 => to_slv(opcode_type, 16#10#),
      844 => to_slv(opcode_type, 16#0A#),
      845 => to_slv(opcode_type, 16#08#),
      846 => to_slv(opcode_type, 16#07#),
      847 => to_slv(opcode_type, 16#06#),
      848 => to_slv(opcode_type, 16#11#),
      849 => to_slv(opcode_type, 16#0C#),
      850 => to_slv(opcode_type, 16#06#),
      851 => to_slv(opcode_type, 16#0B#),
      852 => to_slv(opcode_type, 16#10#),
      853 => to_slv(opcode_type, 16#07#),
      854 => to_slv(opcode_type, 16#08#),
      855 => to_slv(opcode_type, 16#10#),
      856 => to_slv(opcode_type, 16#0B#),
      857 => to_slv(opcode_type, 16#08#),
      858 => to_slv(opcode_type, 16#AE#),
      859 => to_slv(opcode_type, 16#0D#),
      860 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#06#),
      865 => to_slv(opcode_type, 16#08#),
      866 => to_slv(opcode_type, 16#04#),
      867 => to_slv(opcode_type, 16#08#),
      868 => to_slv(opcode_type, 16#0B#),
      869 => to_slv(opcode_type, 16#0D#),
      870 => to_slv(opcode_type, 16#09#),
      871 => to_slv(opcode_type, 16#07#),
      872 => to_slv(opcode_type, 16#EB#),
      873 => to_slv(opcode_type, 16#0B#),
      874 => to_slv(opcode_type, 16#08#),
      875 => to_slv(opcode_type, 16#0F#),
      876 => to_slv(opcode_type, 16#11#),
      877 => to_slv(opcode_type, 16#09#),
      878 => to_slv(opcode_type, 16#08#),
      879 => to_slv(opcode_type, 16#06#),
      880 => to_slv(opcode_type, 16#0F#),
      881 => to_slv(opcode_type, 16#10#),
      882 => to_slv(opcode_type, 16#06#),
      883 => to_slv(opcode_type, 16#0A#),
      884 => to_slv(opcode_type, 16#0D#),
      885 => to_slv(opcode_type, 16#06#),
      886 => to_slv(opcode_type, 16#09#),
      887 => to_slv(opcode_type, 16#11#),
      888 => to_slv(opcode_type, 16#0D#),
      889 => to_slv(opcode_type, 16#09#),
      890 => to_slv(opcode_type, 16#0E#),
      891 => to_slv(opcode_type, 16#10#),
      892 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#07#),
      898 => to_slv(opcode_type, 16#06#),
      899 => to_slv(opcode_type, 16#04#),
      900 => to_slv(opcode_type, 16#0D#),
      901 => to_slv(opcode_type, 16#05#),
      902 => to_slv(opcode_type, 16#0A#),
      903 => to_slv(opcode_type, 16#09#),
      904 => to_slv(opcode_type, 16#09#),
      905 => to_slv(opcode_type, 16#0C#),
      906 => to_slv(opcode_type, 16#0B#),
      907 => to_slv(opcode_type, 16#04#),
      908 => to_slv(opcode_type, 16#11#),
      909 => to_slv(opcode_type, 16#07#),
      910 => to_slv(opcode_type, 16#08#),
      911 => to_slv(opcode_type, 16#07#),
      912 => to_slv(opcode_type, 16#0D#),
      913 => to_slv(opcode_type, 16#D4#),
      914 => to_slv(opcode_type, 16#07#),
      915 => to_slv(opcode_type, 16#0C#),
      916 => to_slv(opcode_type, 16#0D#),
      917 => to_slv(opcode_type, 16#06#),
      918 => to_slv(opcode_type, 16#06#),
      919 => to_slv(opcode_type, 16#0D#),
      920 => to_slv(opcode_type, 16#0D#),
      921 => to_slv(opcode_type, 16#09#),
      922 => to_slv(opcode_type, 16#8D#),
      923 => to_slv(opcode_type, 16#0C#),
      924 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#06#),
      929 => to_slv(opcode_type, 16#08#),
      930 => to_slv(opcode_type, 16#04#),
      931 => to_slv(opcode_type, 16#06#),
      932 => to_slv(opcode_type, 16#0D#),
      933 => to_slv(opcode_type, 16#B5#),
      934 => to_slv(opcode_type, 16#09#),
      935 => to_slv(opcode_type, 16#07#),
      936 => to_slv(opcode_type, 16#11#),
      937 => to_slv(opcode_type, 16#10#),
      938 => to_slv(opcode_type, 16#08#),
      939 => to_slv(opcode_type, 16#11#),
      940 => to_slv(opcode_type, 16#0D#),
      941 => to_slv(opcode_type, 16#07#),
      942 => to_slv(opcode_type, 16#07#),
      943 => to_slv(opcode_type, 16#09#),
      944 => to_slv(opcode_type, 16#62#),
      945 => to_slv(opcode_type, 16#0D#),
      946 => to_slv(opcode_type, 16#06#),
      947 => to_slv(opcode_type, 16#DC#),
      948 => to_slv(opcode_type, 16#0F#),
      949 => to_slv(opcode_type, 16#08#),
      950 => to_slv(opcode_type, 16#06#),
      951 => to_slv(opcode_type, 16#10#),
      952 => to_slv(opcode_type, 16#0A#),
      953 => to_slv(opcode_type, 16#09#),
      954 => to_slv(opcode_type, 16#0D#),
      955 => to_slv(opcode_type, 16#0C#),
      956 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#08#),
      962 => to_slv(opcode_type, 16#03#),
      963 => to_slv(opcode_type, 16#06#),
      964 => to_slv(opcode_type, 16#7B#),
      965 => to_slv(opcode_type, 16#0D#),
      966 => to_slv(opcode_type, 16#06#),
      967 => to_slv(opcode_type, 16#09#),
      968 => to_slv(opcode_type, 16#0C#),
      969 => to_slv(opcode_type, 16#C6#),
      970 => to_slv(opcode_type, 16#08#),
      971 => to_slv(opcode_type, 16#0C#),
      972 => to_slv(opcode_type, 16#6F#),
      973 => to_slv(opcode_type, 16#09#),
      974 => to_slv(opcode_type, 16#08#),
      975 => to_slv(opcode_type, 16#09#),
      976 => to_slv(opcode_type, 16#0B#),
      977 => to_slv(opcode_type, 16#0C#),
      978 => to_slv(opcode_type, 16#09#),
      979 => to_slv(opcode_type, 16#0C#),
      980 => to_slv(opcode_type, 16#0F#),
      981 => to_slv(opcode_type, 16#06#),
      982 => to_slv(opcode_type, 16#09#),
      983 => to_slv(opcode_type, 16#0F#),
      984 => to_slv(opcode_type, 16#0C#),
      985 => to_slv(opcode_type, 16#06#),
      986 => to_slv(opcode_type, 16#0F#),
      987 => to_slv(opcode_type, 16#5C#),
      988 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#06#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#01#),
      995 => to_slv(opcode_type, 16#09#),
      996 => to_slv(opcode_type, 16#11#),
      997 => to_slv(opcode_type, 16#0C#),
      998 => to_slv(opcode_type, 16#07#),
      999 => to_slv(opcode_type, 16#09#),
      1000 => to_slv(opcode_type, 16#0F#),
      1001 => to_slv(opcode_type, 16#0F#),
      1002 => to_slv(opcode_type, 16#06#),
      1003 => to_slv(opcode_type, 16#0C#),
      1004 => to_slv(opcode_type, 16#0F#),
      1005 => to_slv(opcode_type, 16#06#),
      1006 => to_slv(opcode_type, 16#06#),
      1007 => to_slv(opcode_type, 16#06#),
      1008 => to_slv(opcode_type, 16#0E#),
      1009 => to_slv(opcode_type, 16#0B#),
      1010 => to_slv(opcode_type, 16#08#),
      1011 => to_slv(opcode_type, 16#0B#),
      1012 => to_slv(opcode_type, 16#0D#),
      1013 => to_slv(opcode_type, 16#09#),
      1014 => to_slv(opcode_type, 16#06#),
      1015 => to_slv(opcode_type, 16#52#),
      1016 => to_slv(opcode_type, 16#0E#),
      1017 => to_slv(opcode_type, 16#06#),
      1018 => to_slv(opcode_type, 16#11#),
      1019 => to_slv(opcode_type, 16#0F#),
      1020 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#08#),
      1025 => to_slv(opcode_type, 16#08#),
      1026 => to_slv(opcode_type, 16#09#),
      1027 => to_slv(opcode_type, 16#05#),
      1028 => to_slv(opcode_type, 16#10#),
      1029 => to_slv(opcode_type, 16#05#),
      1030 => to_slv(opcode_type, 16#91#),
      1031 => to_slv(opcode_type, 16#09#),
      1032 => to_slv(opcode_type, 16#08#),
      1033 => to_slv(opcode_type, 16#0F#),
      1034 => to_slv(opcode_type, 16#0A#),
      1035 => to_slv(opcode_type, 16#04#),
      1036 => to_slv(opcode_type, 16#10#),
      1037 => to_slv(opcode_type, 16#09#),
      1038 => to_slv(opcode_type, 16#08#),
      1039 => to_slv(opcode_type, 16#08#),
      1040 => to_slv(opcode_type, 16#0D#),
      1041 => to_slv(opcode_type, 16#0B#),
      1042 => to_slv(opcode_type, 16#06#),
      1043 => to_slv(opcode_type, 16#0A#),
      1044 => to_slv(opcode_type, 16#0A#),
      1045 => to_slv(opcode_type, 16#07#),
      1046 => to_slv(opcode_type, 16#09#),
      1047 => to_slv(opcode_type, 16#0C#),
      1048 => to_slv(opcode_type, 16#0F#),
      1049 => to_slv(opcode_type, 16#07#),
      1050 => to_slv(opcode_type, 16#0B#),
      1051 => to_slv(opcode_type, 16#20#),
      1052 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#09#),
      1057 => to_slv(opcode_type, 16#07#),
      1058 => to_slv(opcode_type, 16#09#),
      1059 => to_slv(opcode_type, 16#06#),
      1060 => to_slv(opcode_type, 16#5C#),
      1061 => to_slv(opcode_type, 16#0C#),
      1062 => to_slv(opcode_type, 16#06#),
      1063 => to_slv(opcode_type, 16#10#),
      1064 => to_slv(opcode_type, 16#0D#),
      1065 => to_slv(opcode_type, 16#04#),
      1066 => to_slv(opcode_type, 16#06#),
      1067 => to_slv(opcode_type, 16#0B#),
      1068 => to_slv(opcode_type, 16#0B#),
      1069 => to_slv(opcode_type, 16#08#),
      1070 => to_slv(opcode_type, 16#08#),
      1071 => to_slv(opcode_type, 16#08#),
      1072 => to_slv(opcode_type, 16#10#),
      1073 => to_slv(opcode_type, 16#0D#),
      1074 => to_slv(opcode_type, 16#06#),
      1075 => to_slv(opcode_type, 16#0D#),
      1076 => to_slv(opcode_type, 16#0F#),
      1077 => to_slv(opcode_type, 16#07#),
      1078 => to_slv(opcode_type, 16#06#),
      1079 => to_slv(opcode_type, 16#EA#),
      1080 => to_slv(opcode_type, 16#0D#),
      1081 => to_slv(opcode_type, 16#09#),
      1082 => to_slv(opcode_type, 16#11#),
      1083 => to_slv(opcode_type, 16#0F#),
      1084 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#09#),
      1089 => to_slv(opcode_type, 16#08#),
      1090 => to_slv(opcode_type, 16#03#),
      1091 => to_slv(opcode_type, 16#06#),
      1092 => to_slv(opcode_type, 16#0F#),
      1093 => to_slv(opcode_type, 16#0D#),
      1094 => to_slv(opcode_type, 16#07#),
      1095 => to_slv(opcode_type, 16#09#),
      1096 => to_slv(opcode_type, 16#0B#),
      1097 => to_slv(opcode_type, 16#0C#),
      1098 => to_slv(opcode_type, 16#06#),
      1099 => to_slv(opcode_type, 16#0C#),
      1100 => to_slv(opcode_type, 16#0D#),
      1101 => to_slv(opcode_type, 16#06#),
      1102 => to_slv(opcode_type, 16#09#),
      1103 => to_slv(opcode_type, 16#09#),
      1104 => to_slv(opcode_type, 16#0A#),
      1105 => to_slv(opcode_type, 16#0D#),
      1106 => to_slv(opcode_type, 16#07#),
      1107 => to_slv(opcode_type, 16#11#),
      1108 => to_slv(opcode_type, 16#11#),
      1109 => to_slv(opcode_type, 16#08#),
      1110 => to_slv(opcode_type, 16#07#),
      1111 => to_slv(opcode_type, 16#0E#),
      1112 => to_slv(opcode_type, 16#11#),
      1113 => to_slv(opcode_type, 16#08#),
      1114 => to_slv(opcode_type, 16#10#),
      1115 => to_slv(opcode_type, 16#0C#),
      1116 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#06#),
      1121 => to_slv(opcode_type, 16#09#),
      1122 => to_slv(opcode_type, 16#04#),
      1123 => to_slv(opcode_type, 16#06#),
      1124 => to_slv(opcode_type, 16#CD#),
      1125 => to_slv(opcode_type, 16#10#),
      1126 => to_slv(opcode_type, 16#06#),
      1127 => to_slv(opcode_type, 16#06#),
      1128 => to_slv(opcode_type, 16#0E#),
      1129 => to_slv(opcode_type, 16#10#),
      1130 => to_slv(opcode_type, 16#06#),
      1131 => to_slv(opcode_type, 16#0D#),
      1132 => to_slv(opcode_type, 16#0A#),
      1133 => to_slv(opcode_type, 16#09#),
      1134 => to_slv(opcode_type, 16#06#),
      1135 => to_slv(opcode_type, 16#08#),
      1136 => to_slv(opcode_type, 16#0B#),
      1137 => to_slv(opcode_type, 16#0D#),
      1138 => to_slv(opcode_type, 16#06#),
      1139 => to_slv(opcode_type, 16#10#),
      1140 => to_slv(opcode_type, 16#0C#),
      1141 => to_slv(opcode_type, 16#08#),
      1142 => to_slv(opcode_type, 16#09#),
      1143 => to_slv(opcode_type, 16#0F#),
      1144 => to_slv(opcode_type, 16#0B#),
      1145 => to_slv(opcode_type, 16#08#),
      1146 => to_slv(opcode_type, 16#0C#),
      1147 => to_slv(opcode_type, 16#0F#),
      1148 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#07#),
      1153 => to_slv(opcode_type, 16#09#),
      1154 => to_slv(opcode_type, 16#06#),
      1155 => to_slv(opcode_type, 16#08#),
      1156 => to_slv(opcode_type, 16#C2#),
      1157 => to_slv(opcode_type, 16#0D#),
      1158 => to_slv(opcode_type, 16#04#),
      1159 => to_slv(opcode_type, 16#0A#),
      1160 => to_slv(opcode_type, 16#06#),
      1161 => to_slv(opcode_type, 16#01#),
      1162 => to_slv(opcode_type, 16#0C#),
      1163 => to_slv(opcode_type, 16#05#),
      1164 => to_slv(opcode_type, 16#0E#),
      1165 => to_slv(opcode_type, 16#09#),
      1166 => to_slv(opcode_type, 16#07#),
      1167 => to_slv(opcode_type, 16#09#),
      1168 => to_slv(opcode_type, 16#10#),
      1169 => to_slv(opcode_type, 16#10#),
      1170 => to_slv(opcode_type, 16#09#),
      1171 => to_slv(opcode_type, 16#10#),
      1172 => to_slv(opcode_type, 16#0A#),
      1173 => to_slv(opcode_type, 16#07#),
      1174 => to_slv(opcode_type, 16#07#),
      1175 => to_slv(opcode_type, 16#0C#),
      1176 => to_slv(opcode_type, 16#0C#),
      1177 => to_slv(opcode_type, 16#09#),
      1178 => to_slv(opcode_type, 16#0C#),
      1179 => to_slv(opcode_type, 16#11#),
      1180 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#08#),
      1185 => to_slv(opcode_type, 16#07#),
      1186 => to_slv(opcode_type, 16#09#),
      1187 => to_slv(opcode_type, 16#02#),
      1188 => to_slv(opcode_type, 16#11#),
      1189 => to_slv(opcode_type, 16#03#),
      1190 => to_slv(opcode_type, 16#0F#),
      1191 => to_slv(opcode_type, 16#06#),
      1192 => to_slv(opcode_type, 16#03#),
      1193 => to_slv(opcode_type, 16#0D#),
      1194 => to_slv(opcode_type, 16#06#),
      1195 => to_slv(opcode_type, 16#0D#),
      1196 => to_slv(opcode_type, 16#0B#),
      1197 => to_slv(opcode_type, 16#08#),
      1198 => to_slv(opcode_type, 16#09#),
      1199 => to_slv(opcode_type, 16#09#),
      1200 => to_slv(opcode_type, 16#0F#),
      1201 => to_slv(opcode_type, 16#D2#),
      1202 => to_slv(opcode_type, 16#08#),
      1203 => to_slv(opcode_type, 16#0C#),
      1204 => to_slv(opcode_type, 16#0B#),
      1205 => to_slv(opcode_type, 16#07#),
      1206 => to_slv(opcode_type, 16#07#),
      1207 => to_slv(opcode_type, 16#43#),
      1208 => to_slv(opcode_type, 16#11#),
      1209 => to_slv(opcode_type, 16#07#),
      1210 => to_slv(opcode_type, 16#11#),
      1211 => to_slv(opcode_type, 16#0C#),
      1212 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#09#),
      1217 => to_slv(opcode_type, 16#08#),
      1218 => to_slv(opcode_type, 16#03#),
      1219 => to_slv(opcode_type, 16#08#),
      1220 => to_slv(opcode_type, 16#0B#),
      1221 => to_slv(opcode_type, 16#10#),
      1222 => to_slv(opcode_type, 16#08#),
      1223 => to_slv(opcode_type, 16#06#),
      1224 => to_slv(opcode_type, 16#10#),
      1225 => to_slv(opcode_type, 16#A8#),
      1226 => to_slv(opcode_type, 16#06#),
      1227 => to_slv(opcode_type, 16#10#),
      1228 => to_slv(opcode_type, 16#0C#),
      1229 => to_slv(opcode_type, 16#07#),
      1230 => to_slv(opcode_type, 16#07#),
      1231 => to_slv(opcode_type, 16#09#),
      1232 => to_slv(opcode_type, 16#0D#),
      1233 => to_slv(opcode_type, 16#10#),
      1234 => to_slv(opcode_type, 16#07#),
      1235 => to_slv(opcode_type, 16#0C#),
      1236 => to_slv(opcode_type, 16#0F#),
      1237 => to_slv(opcode_type, 16#06#),
      1238 => to_slv(opcode_type, 16#07#),
      1239 => to_slv(opcode_type, 16#11#),
      1240 => to_slv(opcode_type, 16#0F#),
      1241 => to_slv(opcode_type, 16#08#),
      1242 => to_slv(opcode_type, 16#0C#),
      1243 => to_slv(opcode_type, 16#10#),
      1244 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#09#),
      1249 => to_slv(opcode_type, 16#07#),
      1250 => to_slv(opcode_type, 16#08#),
      1251 => to_slv(opcode_type, 16#05#),
      1252 => to_slv(opcode_type, 16#0E#),
      1253 => to_slv(opcode_type, 16#05#),
      1254 => to_slv(opcode_type, 16#0F#),
      1255 => to_slv(opcode_type, 16#07#),
      1256 => to_slv(opcode_type, 16#04#),
      1257 => to_slv(opcode_type, 16#0C#),
      1258 => to_slv(opcode_type, 16#06#),
      1259 => to_slv(opcode_type, 16#0A#),
      1260 => to_slv(opcode_type, 16#0A#),
      1261 => to_slv(opcode_type, 16#09#),
      1262 => to_slv(opcode_type, 16#07#),
      1263 => to_slv(opcode_type, 16#06#),
      1264 => to_slv(opcode_type, 16#5D#),
      1265 => to_slv(opcode_type, 16#DD#),
      1266 => to_slv(opcode_type, 16#06#),
      1267 => to_slv(opcode_type, 16#0A#),
      1268 => to_slv(opcode_type, 16#11#),
      1269 => to_slv(opcode_type, 16#06#),
      1270 => to_slv(opcode_type, 16#08#),
      1271 => to_slv(opcode_type, 16#0E#),
      1272 => to_slv(opcode_type, 16#0F#),
      1273 => to_slv(opcode_type, 16#08#),
      1274 => to_slv(opcode_type, 16#C8#),
      1275 => to_slv(opcode_type, 16#11#),
      1276 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#07#),
      1281 => to_slv(opcode_type, 16#06#),
      1282 => to_slv(opcode_type, 16#02#),
      1283 => to_slv(opcode_type, 16#08#),
      1284 => to_slv(opcode_type, 16#F9#),
      1285 => to_slv(opcode_type, 16#0C#),
      1286 => to_slv(opcode_type, 16#07#),
      1287 => to_slv(opcode_type, 16#08#),
      1288 => to_slv(opcode_type, 16#0C#),
      1289 => to_slv(opcode_type, 16#11#),
      1290 => to_slv(opcode_type, 16#07#),
      1291 => to_slv(opcode_type, 16#0B#),
      1292 => to_slv(opcode_type, 16#0E#),
      1293 => to_slv(opcode_type, 16#09#),
      1294 => to_slv(opcode_type, 16#06#),
      1295 => to_slv(opcode_type, 16#06#),
      1296 => to_slv(opcode_type, 16#10#),
      1297 => to_slv(opcode_type, 16#0E#),
      1298 => to_slv(opcode_type, 16#06#),
      1299 => to_slv(opcode_type, 16#0F#),
      1300 => to_slv(opcode_type, 16#0D#),
      1301 => to_slv(opcode_type, 16#06#),
      1302 => to_slv(opcode_type, 16#09#),
      1303 => to_slv(opcode_type, 16#0C#),
      1304 => to_slv(opcode_type, 16#0C#),
      1305 => to_slv(opcode_type, 16#06#),
      1306 => to_slv(opcode_type, 16#90#),
      1307 => to_slv(opcode_type, 16#0D#),
      1308 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#08#),
      1313 => to_slv(opcode_type, 16#07#),
      1314 => to_slv(opcode_type, 16#08#),
      1315 => to_slv(opcode_type, 16#08#),
      1316 => to_slv(opcode_type, 16#41#),
      1317 => to_slv(opcode_type, 16#10#),
      1318 => to_slv(opcode_type, 16#06#),
      1319 => to_slv(opcode_type, 16#0D#),
      1320 => to_slv(opcode_type, 16#0C#),
      1321 => to_slv(opcode_type, 16#04#),
      1322 => to_slv(opcode_type, 16#08#),
      1323 => to_slv(opcode_type, 16#0F#),
      1324 => to_slv(opcode_type, 16#11#),
      1325 => to_slv(opcode_type, 16#07#),
      1326 => to_slv(opcode_type, 16#09#),
      1327 => to_slv(opcode_type, 16#07#),
      1328 => to_slv(opcode_type, 16#0D#),
      1329 => to_slv(opcode_type, 16#10#),
      1330 => to_slv(opcode_type, 16#09#),
      1331 => to_slv(opcode_type, 16#E6#),
      1332 => to_slv(opcode_type, 16#0F#),
      1333 => to_slv(opcode_type, 16#07#),
      1334 => to_slv(opcode_type, 16#06#),
      1335 => to_slv(opcode_type, 16#0D#),
      1336 => to_slv(opcode_type, 16#0C#),
      1337 => to_slv(opcode_type, 16#08#),
      1338 => to_slv(opcode_type, 16#0B#),
      1339 => to_slv(opcode_type, 16#0D#),
      1340 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#06#),
      1345 => to_slv(opcode_type, 16#07#),
      1346 => to_slv(opcode_type, 16#08#),
      1347 => to_slv(opcode_type, 16#01#),
      1348 => to_slv(opcode_type, 16#0F#),
      1349 => to_slv(opcode_type, 16#04#),
      1350 => to_slv(opcode_type, 16#0A#),
      1351 => to_slv(opcode_type, 16#06#),
      1352 => to_slv(opcode_type, 16#08#),
      1353 => to_slv(opcode_type, 16#0A#),
      1354 => to_slv(opcode_type, 16#0F#),
      1355 => to_slv(opcode_type, 16#05#),
      1356 => to_slv(opcode_type, 16#CB#),
      1357 => to_slv(opcode_type, 16#09#),
      1358 => to_slv(opcode_type, 16#08#),
      1359 => to_slv(opcode_type, 16#09#),
      1360 => to_slv(opcode_type, 16#11#),
      1361 => to_slv(opcode_type, 16#0B#),
      1362 => to_slv(opcode_type, 16#06#),
      1363 => to_slv(opcode_type, 16#B4#),
      1364 => to_slv(opcode_type, 16#0C#),
      1365 => to_slv(opcode_type, 16#08#),
      1366 => to_slv(opcode_type, 16#09#),
      1367 => to_slv(opcode_type, 16#0D#),
      1368 => to_slv(opcode_type, 16#11#),
      1369 => to_slv(opcode_type, 16#09#),
      1370 => to_slv(opcode_type, 16#0B#),
      1371 => to_slv(opcode_type, 16#0C#),
      1372 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#06#),
      1377 => to_slv(opcode_type, 16#08#),
      1378 => to_slv(opcode_type, 16#01#),
      1379 => to_slv(opcode_type, 16#06#),
      1380 => to_slv(opcode_type, 16#0E#),
      1381 => to_slv(opcode_type, 16#0A#),
      1382 => to_slv(opcode_type, 16#09#),
      1383 => to_slv(opcode_type, 16#06#),
      1384 => to_slv(opcode_type, 16#0A#),
      1385 => to_slv(opcode_type, 16#EC#),
      1386 => to_slv(opcode_type, 16#06#),
      1387 => to_slv(opcode_type, 16#0B#),
      1388 => to_slv(opcode_type, 16#0D#),
      1389 => to_slv(opcode_type, 16#09#),
      1390 => to_slv(opcode_type, 16#08#),
      1391 => to_slv(opcode_type, 16#06#),
      1392 => to_slv(opcode_type, 16#0F#),
      1393 => to_slv(opcode_type, 16#0C#),
      1394 => to_slv(opcode_type, 16#09#),
      1395 => to_slv(opcode_type, 16#B0#),
      1396 => to_slv(opcode_type, 16#0E#),
      1397 => to_slv(opcode_type, 16#09#),
      1398 => to_slv(opcode_type, 16#07#),
      1399 => to_slv(opcode_type, 16#0C#),
      1400 => to_slv(opcode_type, 16#0F#),
      1401 => to_slv(opcode_type, 16#09#),
      1402 => to_slv(opcode_type, 16#0B#),
      1403 => to_slv(opcode_type, 16#0E#),
      1404 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#08#),
      1409 => to_slv(opcode_type, 16#07#),
      1410 => to_slv(opcode_type, 16#09#),
      1411 => to_slv(opcode_type, 16#06#),
      1412 => to_slv(opcode_type, 16#0A#),
      1413 => to_slv(opcode_type, 16#0D#),
      1414 => to_slv(opcode_type, 16#05#),
      1415 => to_slv(opcode_type, 16#10#),
      1416 => to_slv(opcode_type, 16#07#),
      1417 => to_slv(opcode_type, 16#02#),
      1418 => to_slv(opcode_type, 16#93#),
      1419 => to_slv(opcode_type, 16#05#),
      1420 => to_slv(opcode_type, 16#10#),
      1421 => to_slv(opcode_type, 16#06#),
      1422 => to_slv(opcode_type, 16#09#),
      1423 => to_slv(opcode_type, 16#06#),
      1424 => to_slv(opcode_type, 16#0B#),
      1425 => to_slv(opcode_type, 16#0F#),
      1426 => to_slv(opcode_type, 16#09#),
      1427 => to_slv(opcode_type, 16#0B#),
      1428 => to_slv(opcode_type, 16#49#),
      1429 => to_slv(opcode_type, 16#06#),
      1430 => to_slv(opcode_type, 16#09#),
      1431 => to_slv(opcode_type, 16#0A#),
      1432 => to_slv(opcode_type, 16#11#),
      1433 => to_slv(opcode_type, 16#07#),
      1434 => to_slv(opcode_type, 16#0E#),
      1435 => to_slv(opcode_type, 16#81#),
      1436 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#09#),
      1441 => to_slv(opcode_type, 16#07#),
      1442 => to_slv(opcode_type, 16#03#),
      1443 => to_slv(opcode_type, 16#06#),
      1444 => to_slv(opcode_type, 16#6D#),
      1445 => to_slv(opcode_type, 16#0F#),
      1446 => to_slv(opcode_type, 16#09#),
      1447 => to_slv(opcode_type, 16#08#),
      1448 => to_slv(opcode_type, 16#0A#),
      1449 => to_slv(opcode_type, 16#11#),
      1450 => to_slv(opcode_type, 16#09#),
      1451 => to_slv(opcode_type, 16#0E#),
      1452 => to_slv(opcode_type, 16#0B#),
      1453 => to_slv(opcode_type, 16#07#),
      1454 => to_slv(opcode_type, 16#08#),
      1455 => to_slv(opcode_type, 16#09#),
      1456 => to_slv(opcode_type, 16#0B#),
      1457 => to_slv(opcode_type, 16#0F#),
      1458 => to_slv(opcode_type, 16#09#),
      1459 => to_slv(opcode_type, 16#9C#),
      1460 => to_slv(opcode_type, 16#10#),
      1461 => to_slv(opcode_type, 16#09#),
      1462 => to_slv(opcode_type, 16#08#),
      1463 => to_slv(opcode_type, 16#11#),
      1464 => to_slv(opcode_type, 16#0F#),
      1465 => to_slv(opcode_type, 16#08#),
      1466 => to_slv(opcode_type, 16#0C#),
      1467 => to_slv(opcode_type, 16#2B#),
      1468 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#07#),
      1473 => to_slv(opcode_type, 16#09#),
      1474 => to_slv(opcode_type, 16#06#),
      1475 => to_slv(opcode_type, 16#03#),
      1476 => to_slv(opcode_type, 16#0D#),
      1477 => to_slv(opcode_type, 16#04#),
      1478 => to_slv(opcode_type, 16#0D#),
      1479 => to_slv(opcode_type, 16#07#),
      1480 => to_slv(opcode_type, 16#08#),
      1481 => to_slv(opcode_type, 16#1B#),
      1482 => to_slv(opcode_type, 16#0D#),
      1483 => to_slv(opcode_type, 16#06#),
      1484 => to_slv(opcode_type, 16#0B#),
      1485 => to_slv(opcode_type, 16#0A#),
      1486 => to_slv(opcode_type, 16#07#),
      1487 => to_slv(opcode_type, 16#07#),
      1488 => to_slv(opcode_type, 16#09#),
      1489 => to_slv(opcode_type, 16#10#),
      1490 => to_slv(opcode_type, 16#0E#),
      1491 => to_slv(opcode_type, 16#08#),
      1492 => to_slv(opcode_type, 16#0A#),
      1493 => to_slv(opcode_type, 16#0C#),
      1494 => to_slv(opcode_type, 16#07#),
      1495 => to_slv(opcode_type, 16#08#),
      1496 => to_slv(opcode_type, 16#0E#),
      1497 => to_slv(opcode_type, 16#0A#),
      1498 => to_slv(opcode_type, 16#05#),
      1499 => to_slv(opcode_type, 16#0B#),
      1500 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#08#),
      1505 => to_slv(opcode_type, 16#09#),
      1506 => to_slv(opcode_type, 16#07#),
      1507 => to_slv(opcode_type, 16#06#),
      1508 => to_slv(opcode_type, 16#0B#),
      1509 => to_slv(opcode_type, 16#0E#),
      1510 => to_slv(opcode_type, 16#03#),
      1511 => to_slv(opcode_type, 16#0A#),
      1512 => to_slv(opcode_type, 16#08#),
      1513 => to_slv(opcode_type, 16#04#),
      1514 => to_slv(opcode_type, 16#0D#),
      1515 => to_slv(opcode_type, 16#03#),
      1516 => to_slv(opcode_type, 16#0E#),
      1517 => to_slv(opcode_type, 16#08#),
      1518 => to_slv(opcode_type, 16#08#),
      1519 => to_slv(opcode_type, 16#08#),
      1520 => to_slv(opcode_type, 16#0E#),
      1521 => to_slv(opcode_type, 16#0F#),
      1522 => to_slv(opcode_type, 16#07#),
      1523 => to_slv(opcode_type, 16#0D#),
      1524 => to_slv(opcode_type, 16#0D#),
      1525 => to_slv(opcode_type, 16#06#),
      1526 => to_slv(opcode_type, 16#07#),
      1527 => to_slv(opcode_type, 16#0A#),
      1528 => to_slv(opcode_type, 16#0E#),
      1529 => to_slv(opcode_type, 16#07#),
      1530 => to_slv(opcode_type, 16#3E#),
      1531 => to_slv(opcode_type, 16#11#),
      1532 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#06#),
      1537 => to_slv(opcode_type, 16#09#),
      1538 => to_slv(opcode_type, 16#04#),
      1539 => to_slv(opcode_type, 16#07#),
      1540 => to_slv(opcode_type, 16#0B#),
      1541 => to_slv(opcode_type, 16#0D#),
      1542 => to_slv(opcode_type, 16#06#),
      1543 => to_slv(opcode_type, 16#07#),
      1544 => to_slv(opcode_type, 16#0B#),
      1545 => to_slv(opcode_type, 16#0F#),
      1546 => to_slv(opcode_type, 16#06#),
      1547 => to_slv(opcode_type, 16#0B#),
      1548 => to_slv(opcode_type, 16#0C#),
      1549 => to_slv(opcode_type, 16#08#),
      1550 => to_slv(opcode_type, 16#09#),
      1551 => to_slv(opcode_type, 16#09#),
      1552 => to_slv(opcode_type, 16#0B#),
      1553 => to_slv(opcode_type, 16#0E#),
      1554 => to_slv(opcode_type, 16#07#),
      1555 => to_slv(opcode_type, 16#10#),
      1556 => to_slv(opcode_type, 16#0D#),
      1557 => to_slv(opcode_type, 16#06#),
      1558 => to_slv(opcode_type, 16#08#),
      1559 => to_slv(opcode_type, 16#84#),
      1560 => to_slv(opcode_type, 16#0A#),
      1561 => to_slv(opcode_type, 16#08#),
      1562 => to_slv(opcode_type, 16#0D#),
      1563 => to_slv(opcode_type, 16#10#),
      1564 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#08#),
      1569 => to_slv(opcode_type, 16#09#),
      1570 => to_slv(opcode_type, 16#06#),
      1571 => to_slv(opcode_type, 16#06#),
      1572 => to_slv(opcode_type, 16#0C#),
      1573 => to_slv(opcode_type, 16#0E#),
      1574 => to_slv(opcode_type, 16#07#),
      1575 => to_slv(opcode_type, 16#0E#),
      1576 => to_slv(opcode_type, 16#0F#),
      1577 => to_slv(opcode_type, 16#03#),
      1578 => to_slv(opcode_type, 16#06#),
      1579 => to_slv(opcode_type, 16#0C#),
      1580 => to_slv(opcode_type, 16#11#),
      1581 => to_slv(opcode_type, 16#07#),
      1582 => to_slv(opcode_type, 16#07#),
      1583 => to_slv(opcode_type, 16#09#),
      1584 => to_slv(opcode_type, 16#0E#),
      1585 => to_slv(opcode_type, 16#D5#),
      1586 => to_slv(opcode_type, 16#07#),
      1587 => to_slv(opcode_type, 16#11#),
      1588 => to_slv(opcode_type, 16#11#),
      1589 => to_slv(opcode_type, 16#06#),
      1590 => to_slv(opcode_type, 16#08#),
      1591 => to_slv(opcode_type, 16#7B#),
      1592 => to_slv(opcode_type, 16#D7#),
      1593 => to_slv(opcode_type, 16#06#),
      1594 => to_slv(opcode_type, 16#0F#),
      1595 => to_slv(opcode_type, 16#E1#),
      1596 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#07#),
      1602 => to_slv(opcode_type, 16#03#),
      1603 => to_slv(opcode_type, 16#09#),
      1604 => to_slv(opcode_type, 16#0C#),
      1605 => to_slv(opcode_type, 16#0B#),
      1606 => to_slv(opcode_type, 16#06#),
      1607 => to_slv(opcode_type, 16#06#),
      1608 => to_slv(opcode_type, 16#0B#),
      1609 => to_slv(opcode_type, 16#10#),
      1610 => to_slv(opcode_type, 16#09#),
      1611 => to_slv(opcode_type, 16#0F#),
      1612 => to_slv(opcode_type, 16#0E#),
      1613 => to_slv(opcode_type, 16#07#),
      1614 => to_slv(opcode_type, 16#07#),
      1615 => to_slv(opcode_type, 16#09#),
      1616 => to_slv(opcode_type, 16#0D#),
      1617 => to_slv(opcode_type, 16#0E#),
      1618 => to_slv(opcode_type, 16#09#),
      1619 => to_slv(opcode_type, 16#0C#),
      1620 => to_slv(opcode_type, 16#0D#),
      1621 => to_slv(opcode_type, 16#08#),
      1622 => to_slv(opcode_type, 16#06#),
      1623 => to_slv(opcode_type, 16#0C#),
      1624 => to_slv(opcode_type, 16#0A#),
      1625 => to_slv(opcode_type, 16#08#),
      1626 => to_slv(opcode_type, 16#11#),
      1627 => to_slv(opcode_type, 16#0F#),
      1628 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#07#),
      1633 => to_slv(opcode_type, 16#06#),
      1634 => to_slv(opcode_type, 16#08#),
      1635 => to_slv(opcode_type, 16#04#),
      1636 => to_slv(opcode_type, 16#0D#),
      1637 => to_slv(opcode_type, 16#08#),
      1638 => to_slv(opcode_type, 16#0E#),
      1639 => to_slv(opcode_type, 16#C2#),
      1640 => to_slv(opcode_type, 16#07#),
      1641 => to_slv(opcode_type, 16#06#),
      1642 => to_slv(opcode_type, 16#0D#),
      1643 => to_slv(opcode_type, 16#10#),
      1644 => to_slv(opcode_type, 16#05#),
      1645 => to_slv(opcode_type, 16#0B#),
      1646 => to_slv(opcode_type, 16#07#),
      1647 => to_slv(opcode_type, 16#08#),
      1648 => to_slv(opcode_type, 16#03#),
      1649 => to_slv(opcode_type, 16#0B#),
      1650 => to_slv(opcode_type, 16#07#),
      1651 => to_slv(opcode_type, 16#0B#),
      1652 => to_slv(opcode_type, 16#0B#),
      1653 => to_slv(opcode_type, 16#07#),
      1654 => to_slv(opcode_type, 16#06#),
      1655 => to_slv(opcode_type, 16#0B#),
      1656 => to_slv(opcode_type, 16#0E#),
      1657 => to_slv(opcode_type, 16#06#),
      1658 => to_slv(opcode_type, 16#0F#),
      1659 => to_slv(opcode_type, 16#0B#),
      1660 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#09#),
      1666 => to_slv(opcode_type, 16#07#),
      1667 => to_slv(opcode_type, 16#09#),
      1668 => to_slv(opcode_type, 16#0A#),
      1669 => to_slv(opcode_type, 16#0F#),
      1670 => to_slv(opcode_type, 16#09#),
      1671 => to_slv(opcode_type, 16#0A#),
      1672 => to_slv(opcode_type, 16#0D#),
      1673 => to_slv(opcode_type, 16#05#),
      1674 => to_slv(opcode_type, 16#08#),
      1675 => to_slv(opcode_type, 16#10#),
      1676 => to_slv(opcode_type, 16#0D#),
      1677 => to_slv(opcode_type, 16#06#),
      1678 => to_slv(opcode_type, 16#09#),
      1679 => to_slv(opcode_type, 16#07#),
      1680 => to_slv(opcode_type, 16#0C#),
      1681 => to_slv(opcode_type, 16#10#),
      1682 => to_slv(opcode_type, 16#07#),
      1683 => to_slv(opcode_type, 16#5E#),
      1684 => to_slv(opcode_type, 16#0F#),
      1685 => to_slv(opcode_type, 16#06#),
      1686 => to_slv(opcode_type, 16#07#),
      1687 => to_slv(opcode_type, 16#0B#),
      1688 => to_slv(opcode_type, 16#0B#),
      1689 => to_slv(opcode_type, 16#07#),
      1690 => to_slv(opcode_type, 16#F0#),
      1691 => to_slv(opcode_type, 16#0B#),
      1692 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#09#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#05#),
      1699 => to_slv(opcode_type, 16#06#),
      1700 => to_slv(opcode_type, 16#E5#),
      1701 => to_slv(opcode_type, 16#0E#),
      1702 => to_slv(opcode_type, 16#06#),
      1703 => to_slv(opcode_type, 16#09#),
      1704 => to_slv(opcode_type, 16#0E#),
      1705 => to_slv(opcode_type, 16#0F#),
      1706 => to_slv(opcode_type, 16#06#),
      1707 => to_slv(opcode_type, 16#0D#),
      1708 => to_slv(opcode_type, 16#0F#),
      1709 => to_slv(opcode_type, 16#06#),
      1710 => to_slv(opcode_type, 16#06#),
      1711 => to_slv(opcode_type, 16#09#),
      1712 => to_slv(opcode_type, 16#0C#),
      1713 => to_slv(opcode_type, 16#11#),
      1714 => to_slv(opcode_type, 16#09#),
      1715 => to_slv(opcode_type, 16#0F#),
      1716 => to_slv(opcode_type, 16#0F#),
      1717 => to_slv(opcode_type, 16#06#),
      1718 => to_slv(opcode_type, 16#07#),
      1719 => to_slv(opcode_type, 16#0E#),
      1720 => to_slv(opcode_type, 16#0A#),
      1721 => to_slv(opcode_type, 16#07#),
      1722 => to_slv(opcode_type, 16#0C#),
      1723 => to_slv(opcode_type, 16#0F#),
      1724 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#06#),
      1729 => to_slv(opcode_type, 16#07#),
      1730 => to_slv(opcode_type, 16#07#),
      1731 => to_slv(opcode_type, 16#06#),
      1732 => to_slv(opcode_type, 16#0B#),
      1733 => to_slv(opcode_type, 16#F8#),
      1734 => to_slv(opcode_type, 16#02#),
      1735 => to_slv(opcode_type, 16#11#),
      1736 => to_slv(opcode_type, 16#07#),
      1737 => to_slv(opcode_type, 16#03#),
      1738 => to_slv(opcode_type, 16#84#),
      1739 => to_slv(opcode_type, 16#06#),
      1740 => to_slv(opcode_type, 16#10#),
      1741 => to_slv(opcode_type, 16#0D#),
      1742 => to_slv(opcode_type, 16#09#),
      1743 => to_slv(opcode_type, 16#06#),
      1744 => to_slv(opcode_type, 16#05#),
      1745 => to_slv(opcode_type, 16#0C#),
      1746 => to_slv(opcode_type, 16#07#),
      1747 => to_slv(opcode_type, 16#0A#),
      1748 => to_slv(opcode_type, 16#0D#),
      1749 => to_slv(opcode_type, 16#09#),
      1750 => to_slv(opcode_type, 16#07#),
      1751 => to_slv(opcode_type, 16#10#),
      1752 => to_slv(opcode_type, 16#0D#),
      1753 => to_slv(opcode_type, 16#08#),
      1754 => to_slv(opcode_type, 16#0F#),
      1755 => to_slv(opcode_type, 16#0A#),
      1756 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#09#),
      1761 => to_slv(opcode_type, 16#06#),
      1762 => to_slv(opcode_type, 16#01#),
      1763 => to_slv(opcode_type, 16#09#),
      1764 => to_slv(opcode_type, 16#0F#),
      1765 => to_slv(opcode_type, 16#0C#),
      1766 => to_slv(opcode_type, 16#07#),
      1767 => to_slv(opcode_type, 16#09#),
      1768 => to_slv(opcode_type, 16#0A#),
      1769 => to_slv(opcode_type, 16#0C#),
      1770 => to_slv(opcode_type, 16#06#),
      1771 => to_slv(opcode_type, 16#11#),
      1772 => to_slv(opcode_type, 16#0D#),
      1773 => to_slv(opcode_type, 16#06#),
      1774 => to_slv(opcode_type, 16#08#),
      1775 => to_slv(opcode_type, 16#09#),
      1776 => to_slv(opcode_type, 16#0C#),
      1777 => to_slv(opcode_type, 16#0E#),
      1778 => to_slv(opcode_type, 16#08#),
      1779 => to_slv(opcode_type, 16#11#),
      1780 => to_slv(opcode_type, 16#98#),
      1781 => to_slv(opcode_type, 16#07#),
      1782 => to_slv(opcode_type, 16#06#),
      1783 => to_slv(opcode_type, 16#0D#),
      1784 => to_slv(opcode_type, 16#0F#),
      1785 => to_slv(opcode_type, 16#07#),
      1786 => to_slv(opcode_type, 16#0D#),
      1787 => to_slv(opcode_type, 16#10#),
      1788 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#09#),
      1793 => to_slv(opcode_type, 16#08#),
      1794 => to_slv(opcode_type, 16#06#),
      1795 => to_slv(opcode_type, 16#03#),
      1796 => to_slv(opcode_type, 16#10#),
      1797 => to_slv(opcode_type, 16#08#),
      1798 => to_slv(opcode_type, 16#0D#),
      1799 => to_slv(opcode_type, 16#0A#),
      1800 => to_slv(opcode_type, 16#08#),
      1801 => to_slv(opcode_type, 16#06#),
      1802 => to_slv(opcode_type, 16#0B#),
      1803 => to_slv(opcode_type, 16#0D#),
      1804 => to_slv(opcode_type, 16#09#),
      1805 => to_slv(opcode_type, 16#0B#),
      1806 => to_slv(opcode_type, 16#0E#),
      1807 => to_slv(opcode_type, 16#09#),
      1808 => to_slv(opcode_type, 16#06#),
      1809 => to_slv(opcode_type, 16#08#),
      1810 => to_slv(opcode_type, 16#0A#),
      1811 => to_slv(opcode_type, 16#0F#),
      1812 => to_slv(opcode_type, 16#04#),
      1813 => to_slv(opcode_type, 16#10#),
      1814 => to_slv(opcode_type, 16#06#),
      1815 => to_slv(opcode_type, 16#09#),
      1816 => to_slv(opcode_type, 16#79#),
      1817 => to_slv(opcode_type, 16#0B#),
      1818 => to_slv(opcode_type, 16#03#),
      1819 => to_slv(opcode_type, 16#FD#),
      1820 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#09#),
      1825 => to_slv(opcode_type, 16#09#),
      1826 => to_slv(opcode_type, 16#06#),
      1827 => to_slv(opcode_type, 16#06#),
      1828 => to_slv(opcode_type, 16#0D#),
      1829 => to_slv(opcode_type, 16#0F#),
      1830 => to_slv(opcode_type, 16#05#),
      1831 => to_slv(opcode_type, 16#0F#),
      1832 => to_slv(opcode_type, 16#08#),
      1833 => to_slv(opcode_type, 16#07#),
      1834 => to_slv(opcode_type, 16#0C#),
      1835 => to_slv(opcode_type, 16#A6#),
      1836 => to_slv(opcode_type, 16#07#),
      1837 => to_slv(opcode_type, 16#0C#),
      1838 => to_slv(opcode_type, 16#0D#),
      1839 => to_slv(opcode_type, 16#08#),
      1840 => to_slv(opcode_type, 16#08#),
      1841 => to_slv(opcode_type, 16#02#),
      1842 => to_slv(opcode_type, 16#0C#),
      1843 => to_slv(opcode_type, 16#06#),
      1844 => to_slv(opcode_type, 16#0A#),
      1845 => to_slv(opcode_type, 16#11#),
      1846 => to_slv(opcode_type, 16#09#),
      1847 => to_slv(opcode_type, 16#01#),
      1848 => to_slv(opcode_type, 16#11#),
      1849 => to_slv(opcode_type, 16#08#),
      1850 => to_slv(opcode_type, 16#10#),
      1851 => to_slv(opcode_type, 16#8F#),
      1852 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#09#),
      1857 => to_slv(opcode_type, 16#09#),
      1858 => to_slv(opcode_type, 16#05#),
      1859 => to_slv(opcode_type, 16#08#),
      1860 => to_slv(opcode_type, 16#10#),
      1861 => to_slv(opcode_type, 16#0A#),
      1862 => to_slv(opcode_type, 16#07#),
      1863 => to_slv(opcode_type, 16#06#),
      1864 => to_slv(opcode_type, 16#11#),
      1865 => to_slv(opcode_type, 16#0A#),
      1866 => to_slv(opcode_type, 16#09#),
      1867 => to_slv(opcode_type, 16#0E#),
      1868 => to_slv(opcode_type, 16#0F#),
      1869 => to_slv(opcode_type, 16#06#),
      1870 => to_slv(opcode_type, 16#07#),
      1871 => to_slv(opcode_type, 16#08#),
      1872 => to_slv(opcode_type, 16#7E#),
      1873 => to_slv(opcode_type, 16#0C#),
      1874 => to_slv(opcode_type, 16#08#),
      1875 => to_slv(opcode_type, 16#0D#),
      1876 => to_slv(opcode_type, 16#0D#),
      1877 => to_slv(opcode_type, 16#07#),
      1878 => to_slv(opcode_type, 16#09#),
      1879 => to_slv(opcode_type, 16#0E#),
      1880 => to_slv(opcode_type, 16#10#),
      1881 => to_slv(opcode_type, 16#06#),
      1882 => to_slv(opcode_type, 16#0F#),
      1883 => to_slv(opcode_type, 16#0A#),
      1884 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#09#),
      1890 => to_slv(opcode_type, 16#06#),
      1891 => to_slv(opcode_type, 16#09#),
      1892 => to_slv(opcode_type, 16#0A#),
      1893 => to_slv(opcode_type, 16#0E#),
      1894 => to_slv(opcode_type, 16#06#),
      1895 => to_slv(opcode_type, 16#0B#),
      1896 => to_slv(opcode_type, 16#11#),
      1897 => to_slv(opcode_type, 16#06#),
      1898 => to_slv(opcode_type, 16#05#),
      1899 => to_slv(opcode_type, 16#0C#),
      1900 => to_slv(opcode_type, 16#06#),
      1901 => to_slv(opcode_type, 16#0C#),
      1902 => to_slv(opcode_type, 16#10#),
      1903 => to_slv(opcode_type, 16#07#),
      1904 => to_slv(opcode_type, 16#08#),
      1905 => to_slv(opcode_type, 16#07#),
      1906 => to_slv(opcode_type, 16#10#),
      1907 => to_slv(opcode_type, 16#35#),
      1908 => to_slv(opcode_type, 16#05#),
      1909 => to_slv(opcode_type, 16#11#),
      1910 => to_slv(opcode_type, 16#09#),
      1911 => to_slv(opcode_type, 16#09#),
      1912 => to_slv(opcode_type, 16#0F#),
      1913 => to_slv(opcode_type, 16#10#),
      1914 => to_slv(opcode_type, 16#05#),
      1915 => to_slv(opcode_type, 16#0E#),
      1916 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#06#),
      1921 => to_slv(opcode_type, 16#06#),
      1922 => to_slv(opcode_type, 16#03#),
      1923 => to_slv(opcode_type, 16#07#),
      1924 => to_slv(opcode_type, 16#10#),
      1925 => to_slv(opcode_type, 16#0E#),
      1926 => to_slv(opcode_type, 16#09#),
      1927 => to_slv(opcode_type, 16#08#),
      1928 => to_slv(opcode_type, 16#10#),
      1929 => to_slv(opcode_type, 16#0E#),
      1930 => to_slv(opcode_type, 16#08#),
      1931 => to_slv(opcode_type, 16#0F#),
      1932 => to_slv(opcode_type, 16#0D#),
      1933 => to_slv(opcode_type, 16#08#),
      1934 => to_slv(opcode_type, 16#06#),
      1935 => to_slv(opcode_type, 16#06#),
      1936 => to_slv(opcode_type, 16#0D#),
      1937 => to_slv(opcode_type, 16#10#),
      1938 => to_slv(opcode_type, 16#08#),
      1939 => to_slv(opcode_type, 16#0C#),
      1940 => to_slv(opcode_type, 16#10#),
      1941 => to_slv(opcode_type, 16#08#),
      1942 => to_slv(opcode_type, 16#06#),
      1943 => to_slv(opcode_type, 16#10#),
      1944 => to_slv(opcode_type, 16#0E#),
      1945 => to_slv(opcode_type, 16#07#),
      1946 => to_slv(opcode_type, 16#0C#),
      1947 => to_slv(opcode_type, 16#0F#),
      1948 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#07#),
      1953 => to_slv(opcode_type, 16#06#),
      1954 => to_slv(opcode_type, 16#01#),
      1955 => to_slv(opcode_type, 16#07#),
      1956 => to_slv(opcode_type, 16#0D#),
      1957 => to_slv(opcode_type, 16#0A#),
      1958 => to_slv(opcode_type, 16#09#),
      1959 => to_slv(opcode_type, 16#08#),
      1960 => to_slv(opcode_type, 16#0B#),
      1961 => to_slv(opcode_type, 16#79#),
      1962 => to_slv(opcode_type, 16#08#),
      1963 => to_slv(opcode_type, 16#0F#),
      1964 => to_slv(opcode_type, 16#0B#),
      1965 => to_slv(opcode_type, 16#06#),
      1966 => to_slv(opcode_type, 16#09#),
      1967 => to_slv(opcode_type, 16#06#),
      1968 => to_slv(opcode_type, 16#0D#),
      1969 => to_slv(opcode_type, 16#E2#),
      1970 => to_slv(opcode_type, 16#06#),
      1971 => to_slv(opcode_type, 16#0F#),
      1972 => to_slv(opcode_type, 16#0F#),
      1973 => to_slv(opcode_type, 16#06#),
      1974 => to_slv(opcode_type, 16#08#),
      1975 => to_slv(opcode_type, 16#10#),
      1976 => to_slv(opcode_type, 16#0E#),
      1977 => to_slv(opcode_type, 16#09#),
      1978 => to_slv(opcode_type, 16#11#),
      1979 => to_slv(opcode_type, 16#0B#),
      1980 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#07#),
      1985 => to_slv(opcode_type, 16#08#),
      1986 => to_slv(opcode_type, 16#05#),
      1987 => to_slv(opcode_type, 16#07#),
      1988 => to_slv(opcode_type, 16#0F#),
      1989 => to_slv(opcode_type, 16#0D#),
      1990 => to_slv(opcode_type, 16#06#),
      1991 => to_slv(opcode_type, 16#07#),
      1992 => to_slv(opcode_type, 16#0E#),
      1993 => to_slv(opcode_type, 16#0A#),
      1994 => to_slv(opcode_type, 16#09#),
      1995 => to_slv(opcode_type, 16#49#),
      1996 => to_slv(opcode_type, 16#0F#),
      1997 => to_slv(opcode_type, 16#06#),
      1998 => to_slv(opcode_type, 16#08#),
      1999 => to_slv(opcode_type, 16#06#),
      2000 => to_slv(opcode_type, 16#0C#),
      2001 => to_slv(opcode_type, 16#0F#),
      2002 => to_slv(opcode_type, 16#09#),
      2003 => to_slv(opcode_type, 16#10#),
      2004 => to_slv(opcode_type, 16#0A#),
      2005 => to_slv(opcode_type, 16#07#),
      2006 => to_slv(opcode_type, 16#09#),
      2007 => to_slv(opcode_type, 16#0A#),
      2008 => to_slv(opcode_type, 16#0E#),
      2009 => to_slv(opcode_type, 16#08#),
      2010 => to_slv(opcode_type, 16#0B#),
      2011 => to_slv(opcode_type, 16#0C#),
      2012 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#06#),
      2017 => to_slv(opcode_type, 16#07#),
      2018 => to_slv(opcode_type, 16#09#),
      2019 => to_slv(opcode_type, 16#04#),
      2020 => to_slv(opcode_type, 16#11#),
      2021 => to_slv(opcode_type, 16#05#),
      2022 => to_slv(opcode_type, 16#11#),
      2023 => to_slv(opcode_type, 16#08#),
      2024 => to_slv(opcode_type, 16#08#),
      2025 => to_slv(opcode_type, 16#11#),
      2026 => to_slv(opcode_type, 16#CF#),
      2027 => to_slv(opcode_type, 16#01#),
      2028 => to_slv(opcode_type, 16#0D#),
      2029 => to_slv(opcode_type, 16#08#),
      2030 => to_slv(opcode_type, 16#07#),
      2031 => to_slv(opcode_type, 16#07#),
      2032 => to_slv(opcode_type, 16#0C#),
      2033 => to_slv(opcode_type, 16#11#),
      2034 => to_slv(opcode_type, 16#08#),
      2035 => to_slv(opcode_type, 16#11#),
      2036 => to_slv(opcode_type, 16#0D#),
      2037 => to_slv(opcode_type, 16#08#),
      2038 => to_slv(opcode_type, 16#08#),
      2039 => to_slv(opcode_type, 16#0C#),
      2040 => to_slv(opcode_type, 16#0B#),
      2041 => to_slv(opcode_type, 16#06#),
      2042 => to_slv(opcode_type, 16#10#),
      2043 => to_slv(opcode_type, 16#0F#),
      2044 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#06#),
      2049 => to_slv(opcode_type, 16#08#),
      2050 => to_slv(opcode_type, 16#03#),
      2051 => to_slv(opcode_type, 16#08#),
      2052 => to_slv(opcode_type, 16#11#),
      2053 => to_slv(opcode_type, 16#0F#),
      2054 => to_slv(opcode_type, 16#07#),
      2055 => to_slv(opcode_type, 16#09#),
      2056 => to_slv(opcode_type, 16#11#),
      2057 => to_slv(opcode_type, 16#0E#),
      2058 => to_slv(opcode_type, 16#09#),
      2059 => to_slv(opcode_type, 16#0B#),
      2060 => to_slv(opcode_type, 16#0A#),
      2061 => to_slv(opcode_type, 16#07#),
      2062 => to_slv(opcode_type, 16#07#),
      2063 => to_slv(opcode_type, 16#06#),
      2064 => to_slv(opcode_type, 16#0F#),
      2065 => to_slv(opcode_type, 16#0C#),
      2066 => to_slv(opcode_type, 16#08#),
      2067 => to_slv(opcode_type, 16#11#),
      2068 => to_slv(opcode_type, 16#0E#),
      2069 => to_slv(opcode_type, 16#07#),
      2070 => to_slv(opcode_type, 16#06#),
      2071 => to_slv(opcode_type, 16#11#),
      2072 => to_slv(opcode_type, 16#0A#),
      2073 => to_slv(opcode_type, 16#08#),
      2074 => to_slv(opcode_type, 16#10#),
      2075 => to_slv(opcode_type, 16#0A#),
      2076 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#08#),
      2081 => to_slv(opcode_type, 16#09#),
      2082 => to_slv(opcode_type, 16#04#),
      2083 => to_slv(opcode_type, 16#07#),
      2084 => to_slv(opcode_type, 16#0B#),
      2085 => to_slv(opcode_type, 16#0C#),
      2086 => to_slv(opcode_type, 16#09#),
      2087 => to_slv(opcode_type, 16#08#),
      2088 => to_slv(opcode_type, 16#0C#),
      2089 => to_slv(opcode_type, 16#0A#),
      2090 => to_slv(opcode_type, 16#08#),
      2091 => to_slv(opcode_type, 16#0B#),
      2092 => to_slv(opcode_type, 16#0C#),
      2093 => to_slv(opcode_type, 16#07#),
      2094 => to_slv(opcode_type, 16#07#),
      2095 => to_slv(opcode_type, 16#07#),
      2096 => to_slv(opcode_type, 16#0D#),
      2097 => to_slv(opcode_type, 16#0D#),
      2098 => to_slv(opcode_type, 16#08#),
      2099 => to_slv(opcode_type, 16#0C#),
      2100 => to_slv(opcode_type, 16#11#),
      2101 => to_slv(opcode_type, 16#06#),
      2102 => to_slv(opcode_type, 16#08#),
      2103 => to_slv(opcode_type, 16#0E#),
      2104 => to_slv(opcode_type, 16#0D#),
      2105 => to_slv(opcode_type, 16#08#),
      2106 => to_slv(opcode_type, 16#0E#),
      2107 => to_slv(opcode_type, 16#0A#),
      2108 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#06#),
      2113 => to_slv(opcode_type, 16#09#),
      2114 => to_slv(opcode_type, 16#05#),
      2115 => to_slv(opcode_type, 16#08#),
      2116 => to_slv(opcode_type, 16#0C#),
      2117 => to_slv(opcode_type, 16#10#),
      2118 => to_slv(opcode_type, 16#07#),
      2119 => to_slv(opcode_type, 16#06#),
      2120 => to_slv(opcode_type, 16#0F#),
      2121 => to_slv(opcode_type, 16#0D#),
      2122 => to_slv(opcode_type, 16#07#),
      2123 => to_slv(opcode_type, 16#0A#),
      2124 => to_slv(opcode_type, 16#0F#),
      2125 => to_slv(opcode_type, 16#09#),
      2126 => to_slv(opcode_type, 16#06#),
      2127 => to_slv(opcode_type, 16#08#),
      2128 => to_slv(opcode_type, 16#0B#),
      2129 => to_slv(opcode_type, 16#0D#),
      2130 => to_slv(opcode_type, 16#08#),
      2131 => to_slv(opcode_type, 16#0C#),
      2132 => to_slv(opcode_type, 16#0E#),
      2133 => to_slv(opcode_type, 16#07#),
      2134 => to_slv(opcode_type, 16#08#),
      2135 => to_slv(opcode_type, 16#11#),
      2136 => to_slv(opcode_type, 16#11#),
      2137 => to_slv(opcode_type, 16#06#),
      2138 => to_slv(opcode_type, 16#0D#),
      2139 => to_slv(opcode_type, 16#0E#),
      2140 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#07#),
      2145 => to_slv(opcode_type, 16#06#),
      2146 => to_slv(opcode_type, 16#07#),
      2147 => to_slv(opcode_type, 16#06#),
      2148 => to_slv(opcode_type, 16#0A#),
      2149 => to_slv(opcode_type, 16#0B#),
      2150 => to_slv(opcode_type, 16#07#),
      2151 => to_slv(opcode_type, 16#0F#),
      2152 => to_slv(opcode_type, 16#0F#),
      2153 => to_slv(opcode_type, 16#07#),
      2154 => to_slv(opcode_type, 16#09#),
      2155 => to_slv(opcode_type, 16#0C#),
      2156 => to_slv(opcode_type, 16#11#),
      2157 => to_slv(opcode_type, 16#08#),
      2158 => to_slv(opcode_type, 16#0A#),
      2159 => to_slv(opcode_type, 16#0D#),
      2160 => to_slv(opcode_type, 16#07#),
      2161 => to_slv(opcode_type, 16#04#),
      2162 => to_slv(opcode_type, 16#09#),
      2163 => to_slv(opcode_type, 16#1F#),
      2164 => to_slv(opcode_type, 16#0C#),
      2165 => to_slv(opcode_type, 16#09#),
      2166 => to_slv(opcode_type, 16#09#),
      2167 => to_slv(opcode_type, 16#10#),
      2168 => to_slv(opcode_type, 16#0F#),
      2169 => to_slv(opcode_type, 16#07#),
      2170 => to_slv(opcode_type, 16#0E#),
      2171 => to_slv(opcode_type, 16#0B#),
      2172 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#09#),
      2177 => to_slv(opcode_type, 16#06#),
      2178 => to_slv(opcode_type, 16#04#),
      2179 => to_slv(opcode_type, 16#06#),
      2180 => to_slv(opcode_type, 16#0C#),
      2181 => to_slv(opcode_type, 16#11#),
      2182 => to_slv(opcode_type, 16#06#),
      2183 => to_slv(opcode_type, 16#07#),
      2184 => to_slv(opcode_type, 16#D0#),
      2185 => to_slv(opcode_type, 16#0F#),
      2186 => to_slv(opcode_type, 16#06#),
      2187 => to_slv(opcode_type, 16#0C#),
      2188 => to_slv(opcode_type, 16#0E#),
      2189 => to_slv(opcode_type, 16#06#),
      2190 => to_slv(opcode_type, 16#08#),
      2191 => to_slv(opcode_type, 16#08#),
      2192 => to_slv(opcode_type, 16#0F#),
      2193 => to_slv(opcode_type, 16#0C#),
      2194 => to_slv(opcode_type, 16#09#),
      2195 => to_slv(opcode_type, 16#A3#),
      2196 => to_slv(opcode_type, 16#10#),
      2197 => to_slv(opcode_type, 16#08#),
      2198 => to_slv(opcode_type, 16#06#),
      2199 => to_slv(opcode_type, 16#0E#),
      2200 => to_slv(opcode_type, 16#0A#),
      2201 => to_slv(opcode_type, 16#07#),
      2202 => to_slv(opcode_type, 16#0C#),
      2203 => to_slv(opcode_type, 16#0A#),
      2204 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#08#),
      2209 => to_slv(opcode_type, 16#09#),
      2210 => to_slv(opcode_type, 16#08#),
      2211 => to_slv(opcode_type, 16#07#),
      2212 => to_slv(opcode_type, 16#0E#),
      2213 => to_slv(opcode_type, 16#0F#),
      2214 => to_slv(opcode_type, 16#08#),
      2215 => to_slv(opcode_type, 16#0F#),
      2216 => to_slv(opcode_type, 16#0E#),
      2217 => to_slv(opcode_type, 16#02#),
      2218 => to_slv(opcode_type, 16#09#),
      2219 => to_slv(opcode_type, 16#0F#),
      2220 => to_slv(opcode_type, 16#10#),
      2221 => to_slv(opcode_type, 16#07#),
      2222 => to_slv(opcode_type, 16#07#),
      2223 => to_slv(opcode_type, 16#07#),
      2224 => to_slv(opcode_type, 16#0C#),
      2225 => to_slv(opcode_type, 16#0D#),
      2226 => to_slv(opcode_type, 16#09#),
      2227 => to_slv(opcode_type, 16#0C#),
      2228 => to_slv(opcode_type, 16#0E#),
      2229 => to_slv(opcode_type, 16#09#),
      2230 => to_slv(opcode_type, 16#07#),
      2231 => to_slv(opcode_type, 16#0B#),
      2232 => to_slv(opcode_type, 16#86#),
      2233 => to_slv(opcode_type, 16#08#),
      2234 => to_slv(opcode_type, 16#0B#),
      2235 => to_slv(opcode_type, 16#B5#),
      2236 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#09#),
      2241 => to_slv(opcode_type, 16#06#),
      2242 => to_slv(opcode_type, 16#06#),
      2243 => to_slv(opcode_type, 16#02#),
      2244 => to_slv(opcode_type, 16#0A#),
      2245 => to_slv(opcode_type, 16#06#),
      2246 => to_slv(opcode_type, 16#0A#),
      2247 => to_slv(opcode_type, 16#0E#),
      2248 => to_slv(opcode_type, 16#09#),
      2249 => to_slv(opcode_type, 16#02#),
      2250 => to_slv(opcode_type, 16#0C#),
      2251 => to_slv(opcode_type, 16#06#),
      2252 => to_slv(opcode_type, 16#0E#),
      2253 => to_slv(opcode_type, 16#10#),
      2254 => to_slv(opcode_type, 16#09#),
      2255 => to_slv(opcode_type, 16#09#),
      2256 => to_slv(opcode_type, 16#07#),
      2257 => to_slv(opcode_type, 16#0A#),
      2258 => to_slv(opcode_type, 16#0D#),
      2259 => to_slv(opcode_type, 16#01#),
      2260 => to_slv(opcode_type, 16#0F#),
      2261 => to_slv(opcode_type, 16#07#),
      2262 => to_slv(opcode_type, 16#07#),
      2263 => to_slv(opcode_type, 16#0C#),
      2264 => to_slv(opcode_type, 16#0F#),
      2265 => to_slv(opcode_type, 16#08#),
      2266 => to_slv(opcode_type, 16#C4#),
      2267 => to_slv(opcode_type, 16#0F#),
      2268 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#07#),
      2273 => to_slv(opcode_type, 16#09#),
      2274 => to_slv(opcode_type, 16#04#),
      2275 => to_slv(opcode_type, 16#06#),
      2276 => to_slv(opcode_type, 16#0A#),
      2277 => to_slv(opcode_type, 16#0E#),
      2278 => to_slv(opcode_type, 16#09#),
      2279 => to_slv(opcode_type, 16#06#),
      2280 => to_slv(opcode_type, 16#0C#),
      2281 => to_slv(opcode_type, 16#0E#),
      2282 => to_slv(opcode_type, 16#08#),
      2283 => to_slv(opcode_type, 16#0C#),
      2284 => to_slv(opcode_type, 16#0C#),
      2285 => to_slv(opcode_type, 16#09#),
      2286 => to_slv(opcode_type, 16#06#),
      2287 => to_slv(opcode_type, 16#08#),
      2288 => to_slv(opcode_type, 16#AB#),
      2289 => to_slv(opcode_type, 16#0F#),
      2290 => to_slv(opcode_type, 16#09#),
      2291 => to_slv(opcode_type, 16#0E#),
      2292 => to_slv(opcode_type, 16#FF#),
      2293 => to_slv(opcode_type, 16#07#),
      2294 => to_slv(opcode_type, 16#09#),
      2295 => to_slv(opcode_type, 16#0D#),
      2296 => to_slv(opcode_type, 16#11#),
      2297 => to_slv(opcode_type, 16#07#),
      2298 => to_slv(opcode_type, 16#0E#),
      2299 => to_slv(opcode_type, 16#10#),
      2300 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#09#),
      2305 => to_slv(opcode_type, 16#09#),
      2306 => to_slv(opcode_type, 16#04#),
      2307 => to_slv(opcode_type, 16#08#),
      2308 => to_slv(opcode_type, 16#0D#),
      2309 => to_slv(opcode_type, 16#10#),
      2310 => to_slv(opcode_type, 16#07#),
      2311 => to_slv(opcode_type, 16#08#),
      2312 => to_slv(opcode_type, 16#10#),
      2313 => to_slv(opcode_type, 16#10#),
      2314 => to_slv(opcode_type, 16#09#),
      2315 => to_slv(opcode_type, 16#11#),
      2316 => to_slv(opcode_type, 16#11#),
      2317 => to_slv(opcode_type, 16#08#),
      2318 => to_slv(opcode_type, 16#09#),
      2319 => to_slv(opcode_type, 16#08#),
      2320 => to_slv(opcode_type, 16#10#),
      2321 => to_slv(opcode_type, 16#0A#),
      2322 => to_slv(opcode_type, 16#06#),
      2323 => to_slv(opcode_type, 16#D8#),
      2324 => to_slv(opcode_type, 16#0B#),
      2325 => to_slv(opcode_type, 16#07#),
      2326 => to_slv(opcode_type, 16#06#),
      2327 => to_slv(opcode_type, 16#0F#),
      2328 => to_slv(opcode_type, 16#0D#),
      2329 => to_slv(opcode_type, 16#07#),
      2330 => to_slv(opcode_type, 16#6F#),
      2331 => to_slv(opcode_type, 16#0F#),
      2332 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#09#),
      2337 => to_slv(opcode_type, 16#07#),
      2338 => to_slv(opcode_type, 16#03#),
      2339 => to_slv(opcode_type, 16#08#),
      2340 => to_slv(opcode_type, 16#11#),
      2341 => to_slv(opcode_type, 16#0D#),
      2342 => to_slv(opcode_type, 16#07#),
      2343 => to_slv(opcode_type, 16#06#),
      2344 => to_slv(opcode_type, 16#10#),
      2345 => to_slv(opcode_type, 16#0A#),
      2346 => to_slv(opcode_type, 16#09#),
      2347 => to_slv(opcode_type, 16#0E#),
      2348 => to_slv(opcode_type, 16#0C#),
      2349 => to_slv(opcode_type, 16#09#),
      2350 => to_slv(opcode_type, 16#09#),
      2351 => to_slv(opcode_type, 16#06#),
      2352 => to_slv(opcode_type, 16#0F#),
      2353 => to_slv(opcode_type, 16#11#),
      2354 => to_slv(opcode_type, 16#09#),
      2355 => to_slv(opcode_type, 16#0A#),
      2356 => to_slv(opcode_type, 16#0F#),
      2357 => to_slv(opcode_type, 16#08#),
      2358 => to_slv(opcode_type, 16#07#),
      2359 => to_slv(opcode_type, 16#0B#),
      2360 => to_slv(opcode_type, 16#0D#),
      2361 => to_slv(opcode_type, 16#07#),
      2362 => to_slv(opcode_type, 16#0C#),
      2363 => to_slv(opcode_type, 16#88#),
      2364 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#07#),
      2369 => to_slv(opcode_type, 16#06#),
      2370 => to_slv(opcode_type, 16#01#),
      2371 => to_slv(opcode_type, 16#09#),
      2372 => to_slv(opcode_type, 16#0D#),
      2373 => to_slv(opcode_type, 16#4F#),
      2374 => to_slv(opcode_type, 16#07#),
      2375 => to_slv(opcode_type, 16#07#),
      2376 => to_slv(opcode_type, 16#0E#),
      2377 => to_slv(opcode_type, 16#0F#),
      2378 => to_slv(opcode_type, 16#08#),
      2379 => to_slv(opcode_type, 16#10#),
      2380 => to_slv(opcode_type, 16#0F#),
      2381 => to_slv(opcode_type, 16#08#),
      2382 => to_slv(opcode_type, 16#06#),
      2383 => to_slv(opcode_type, 16#08#),
      2384 => to_slv(opcode_type, 16#0B#),
      2385 => to_slv(opcode_type, 16#0E#),
      2386 => to_slv(opcode_type, 16#09#),
      2387 => to_slv(opcode_type, 16#5D#),
      2388 => to_slv(opcode_type, 16#0B#),
      2389 => to_slv(opcode_type, 16#06#),
      2390 => to_slv(opcode_type, 16#07#),
      2391 => to_slv(opcode_type, 16#10#),
      2392 => to_slv(opcode_type, 16#11#),
      2393 => to_slv(opcode_type, 16#06#),
      2394 => to_slv(opcode_type, 16#0B#),
      2395 => to_slv(opcode_type, 16#0B#),
      2396 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#07#),
      2402 => to_slv(opcode_type, 16#08#),
      2403 => to_slv(opcode_type, 16#07#),
      2404 => to_slv(opcode_type, 16#0E#),
      2405 => to_slv(opcode_type, 16#0A#),
      2406 => to_slv(opcode_type, 16#08#),
      2407 => to_slv(opcode_type, 16#0F#),
      2408 => to_slv(opcode_type, 16#0A#),
      2409 => to_slv(opcode_type, 16#06#),
      2410 => to_slv(opcode_type, 16#04#),
      2411 => to_slv(opcode_type, 16#0F#),
      2412 => to_slv(opcode_type, 16#05#),
      2413 => to_slv(opcode_type, 16#0C#),
      2414 => to_slv(opcode_type, 16#06#),
      2415 => to_slv(opcode_type, 16#08#),
      2416 => to_slv(opcode_type, 16#02#),
      2417 => to_slv(opcode_type, 16#10#),
      2418 => to_slv(opcode_type, 16#07#),
      2419 => to_slv(opcode_type, 16#0E#),
      2420 => to_slv(opcode_type, 16#0C#),
      2421 => to_slv(opcode_type, 16#08#),
      2422 => to_slv(opcode_type, 16#09#),
      2423 => to_slv(opcode_type, 16#0E#),
      2424 => to_slv(opcode_type, 16#6E#),
      2425 => to_slv(opcode_type, 16#07#),
      2426 => to_slv(opcode_type, 16#10#),
      2427 => to_slv(opcode_type, 16#11#),
      2428 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#08#),
      2433 => to_slv(opcode_type, 16#07#),
      2434 => to_slv(opcode_type, 16#04#),
      2435 => to_slv(opcode_type, 16#06#),
      2436 => to_slv(opcode_type, 16#10#),
      2437 => to_slv(opcode_type, 16#0F#),
      2438 => to_slv(opcode_type, 16#08#),
      2439 => to_slv(opcode_type, 16#07#),
      2440 => to_slv(opcode_type, 16#10#),
      2441 => to_slv(opcode_type, 16#0F#),
      2442 => to_slv(opcode_type, 16#09#),
      2443 => to_slv(opcode_type, 16#0C#),
      2444 => to_slv(opcode_type, 16#0B#),
      2445 => to_slv(opcode_type, 16#07#),
      2446 => to_slv(opcode_type, 16#07#),
      2447 => to_slv(opcode_type, 16#06#),
      2448 => to_slv(opcode_type, 16#11#),
      2449 => to_slv(opcode_type, 16#0E#),
      2450 => to_slv(opcode_type, 16#07#),
      2451 => to_slv(opcode_type, 16#0F#),
      2452 => to_slv(opcode_type, 16#0E#),
      2453 => to_slv(opcode_type, 16#08#),
      2454 => to_slv(opcode_type, 16#08#),
      2455 => to_slv(opcode_type, 16#0B#),
      2456 => to_slv(opcode_type, 16#41#),
      2457 => to_slv(opcode_type, 16#09#),
      2458 => to_slv(opcode_type, 16#0B#),
      2459 => to_slv(opcode_type, 16#0C#),
      2460 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#08#),
      2465 => to_slv(opcode_type, 16#06#),
      2466 => to_slv(opcode_type, 16#07#),
      2467 => to_slv(opcode_type, 16#04#),
      2468 => to_slv(opcode_type, 16#11#),
      2469 => to_slv(opcode_type, 16#04#),
      2470 => to_slv(opcode_type, 16#0E#),
      2471 => to_slv(opcode_type, 16#08#),
      2472 => to_slv(opcode_type, 16#07#),
      2473 => to_slv(opcode_type, 16#11#),
      2474 => to_slv(opcode_type, 16#10#),
      2475 => to_slv(opcode_type, 16#02#),
      2476 => to_slv(opcode_type, 16#0B#),
      2477 => to_slv(opcode_type, 16#07#),
      2478 => to_slv(opcode_type, 16#08#),
      2479 => to_slv(opcode_type, 16#07#),
      2480 => to_slv(opcode_type, 16#0C#),
      2481 => to_slv(opcode_type, 16#11#),
      2482 => to_slv(opcode_type, 16#09#),
      2483 => to_slv(opcode_type, 16#0D#),
      2484 => to_slv(opcode_type, 16#0B#),
      2485 => to_slv(opcode_type, 16#08#),
      2486 => to_slv(opcode_type, 16#08#),
      2487 => to_slv(opcode_type, 16#E8#),
      2488 => to_slv(opcode_type, 16#A5#),
      2489 => to_slv(opcode_type, 16#06#),
      2490 => to_slv(opcode_type, 16#0C#),
      2491 => to_slv(opcode_type, 16#10#),
      2492 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#07#),
      2497 => to_slv(opcode_type, 16#07#),
      2498 => to_slv(opcode_type, 16#01#),
      2499 => to_slv(opcode_type, 16#07#),
      2500 => to_slv(opcode_type, 16#22#),
      2501 => to_slv(opcode_type, 16#0D#),
      2502 => to_slv(opcode_type, 16#08#),
      2503 => to_slv(opcode_type, 16#09#),
      2504 => to_slv(opcode_type, 16#85#),
      2505 => to_slv(opcode_type, 16#11#),
      2506 => to_slv(opcode_type, 16#07#),
      2507 => to_slv(opcode_type, 16#0B#),
      2508 => to_slv(opcode_type, 16#0C#),
      2509 => to_slv(opcode_type, 16#09#),
      2510 => to_slv(opcode_type, 16#06#),
      2511 => to_slv(opcode_type, 16#08#),
      2512 => to_slv(opcode_type, 16#0F#),
      2513 => to_slv(opcode_type, 16#10#),
      2514 => to_slv(opcode_type, 16#08#),
      2515 => to_slv(opcode_type, 16#54#),
      2516 => to_slv(opcode_type, 16#0D#),
      2517 => to_slv(opcode_type, 16#06#),
      2518 => to_slv(opcode_type, 16#06#),
      2519 => to_slv(opcode_type, 16#0D#),
      2520 => to_slv(opcode_type, 16#18#),
      2521 => to_slv(opcode_type, 16#07#),
      2522 => to_slv(opcode_type, 16#0B#),
      2523 => to_slv(opcode_type, 16#30#),
      2524 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#08#),
      2530 => to_slv(opcode_type, 16#02#),
      2531 => to_slv(opcode_type, 16#07#),
      2532 => to_slv(opcode_type, 16#11#),
      2533 => to_slv(opcode_type, 16#88#),
      2534 => to_slv(opcode_type, 16#08#),
      2535 => to_slv(opcode_type, 16#09#),
      2536 => to_slv(opcode_type, 16#0A#),
      2537 => to_slv(opcode_type, 16#0B#),
      2538 => to_slv(opcode_type, 16#09#),
      2539 => to_slv(opcode_type, 16#0D#),
      2540 => to_slv(opcode_type, 16#0B#),
      2541 => to_slv(opcode_type, 16#08#),
      2542 => to_slv(opcode_type, 16#06#),
      2543 => to_slv(opcode_type, 16#07#),
      2544 => to_slv(opcode_type, 16#0F#),
      2545 => to_slv(opcode_type, 16#0E#),
      2546 => to_slv(opcode_type, 16#09#),
      2547 => to_slv(opcode_type, 16#0E#),
      2548 => to_slv(opcode_type, 16#11#),
      2549 => to_slv(opcode_type, 16#09#),
      2550 => to_slv(opcode_type, 16#09#),
      2551 => to_slv(opcode_type, 16#49#),
      2552 => to_slv(opcode_type, 16#0A#),
      2553 => to_slv(opcode_type, 16#08#),
      2554 => to_slv(opcode_type, 16#0B#),
      2555 => to_slv(opcode_type, 16#FB#),
      2556 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#06#),
      2561 => to_slv(opcode_type, 16#06#),
      2562 => to_slv(opcode_type, 16#09#),
      2563 => to_slv(opcode_type, 16#06#),
      2564 => to_slv(opcode_type, 16#0F#),
      2565 => to_slv(opcode_type, 16#0A#),
      2566 => to_slv(opcode_type, 16#07#),
      2567 => to_slv(opcode_type, 16#0D#),
      2568 => to_slv(opcode_type, 16#0A#),
      2569 => to_slv(opcode_type, 16#01#),
      2570 => to_slv(opcode_type, 16#06#),
      2571 => to_slv(opcode_type, 16#0A#),
      2572 => to_slv(opcode_type, 16#11#),
      2573 => to_slv(opcode_type, 16#07#),
      2574 => to_slv(opcode_type, 16#07#),
      2575 => to_slv(opcode_type, 16#08#),
      2576 => to_slv(opcode_type, 16#23#),
      2577 => to_slv(opcode_type, 16#0C#),
      2578 => to_slv(opcode_type, 16#08#),
      2579 => to_slv(opcode_type, 16#35#),
      2580 => to_slv(opcode_type, 16#10#),
      2581 => to_slv(opcode_type, 16#07#),
      2582 => to_slv(opcode_type, 16#06#),
      2583 => to_slv(opcode_type, 16#0B#),
      2584 => to_slv(opcode_type, 16#C2#),
      2585 => to_slv(opcode_type, 16#08#),
      2586 => to_slv(opcode_type, 16#0B#),
      2587 => to_slv(opcode_type, 16#10#),
      2588 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#08#),
      2593 => to_slv(opcode_type, 16#07#),
      2594 => to_slv(opcode_type, 16#05#),
      2595 => to_slv(opcode_type, 16#08#),
      2596 => to_slv(opcode_type, 16#0C#),
      2597 => to_slv(opcode_type, 16#0D#),
      2598 => to_slv(opcode_type, 16#09#),
      2599 => to_slv(opcode_type, 16#06#),
      2600 => to_slv(opcode_type, 16#0C#),
      2601 => to_slv(opcode_type, 16#0F#),
      2602 => to_slv(opcode_type, 16#09#),
      2603 => to_slv(opcode_type, 16#11#),
      2604 => to_slv(opcode_type, 16#0D#),
      2605 => to_slv(opcode_type, 16#07#),
      2606 => to_slv(opcode_type, 16#08#),
      2607 => to_slv(opcode_type, 16#08#),
      2608 => to_slv(opcode_type, 16#0B#),
      2609 => to_slv(opcode_type, 16#82#),
      2610 => to_slv(opcode_type, 16#08#),
      2611 => to_slv(opcode_type, 16#0C#),
      2612 => to_slv(opcode_type, 16#4F#),
      2613 => to_slv(opcode_type, 16#09#),
      2614 => to_slv(opcode_type, 16#08#),
      2615 => to_slv(opcode_type, 16#0E#),
      2616 => to_slv(opcode_type, 16#0E#),
      2617 => to_slv(opcode_type, 16#09#),
      2618 => to_slv(opcode_type, 16#0A#),
      2619 => to_slv(opcode_type, 16#11#),
      2620 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#08#),
      2625 => to_slv(opcode_type, 16#09#),
      2626 => to_slv(opcode_type, 16#08#),
      2627 => to_slv(opcode_type, 16#05#),
      2628 => to_slv(opcode_type, 16#0F#),
      2629 => to_slv(opcode_type, 16#03#),
      2630 => to_slv(opcode_type, 16#0B#),
      2631 => to_slv(opcode_type, 16#07#),
      2632 => to_slv(opcode_type, 16#07#),
      2633 => to_slv(opcode_type, 16#0A#),
      2634 => to_slv(opcode_type, 16#0E#),
      2635 => to_slv(opcode_type, 16#01#),
      2636 => to_slv(opcode_type, 16#D9#),
      2637 => to_slv(opcode_type, 16#09#),
      2638 => to_slv(opcode_type, 16#06#),
      2639 => to_slv(opcode_type, 16#08#),
      2640 => to_slv(opcode_type, 16#0B#),
      2641 => to_slv(opcode_type, 16#0A#),
      2642 => to_slv(opcode_type, 16#07#),
      2643 => to_slv(opcode_type, 16#0F#),
      2644 => to_slv(opcode_type, 16#0B#),
      2645 => to_slv(opcode_type, 16#06#),
      2646 => to_slv(opcode_type, 16#09#),
      2647 => to_slv(opcode_type, 16#0B#),
      2648 => to_slv(opcode_type, 16#0F#),
      2649 => to_slv(opcode_type, 16#09#),
      2650 => to_slv(opcode_type, 16#0A#),
      2651 => to_slv(opcode_type, 16#0B#),
      2652 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#09#),
      2657 => to_slv(opcode_type, 16#08#),
      2658 => to_slv(opcode_type, 16#07#),
      2659 => to_slv(opcode_type, 16#09#),
      2660 => to_slv(opcode_type, 16#10#),
      2661 => to_slv(opcode_type, 16#0F#),
      2662 => to_slv(opcode_type, 16#02#),
      2663 => to_slv(opcode_type, 16#0A#),
      2664 => to_slv(opcode_type, 16#08#),
      2665 => to_slv(opcode_type, 16#06#),
      2666 => to_slv(opcode_type, 16#10#),
      2667 => to_slv(opcode_type, 16#CE#),
      2668 => to_slv(opcode_type, 16#03#),
      2669 => to_slv(opcode_type, 16#0E#),
      2670 => to_slv(opcode_type, 16#07#),
      2671 => to_slv(opcode_type, 16#08#),
      2672 => to_slv(opcode_type, 16#09#),
      2673 => to_slv(opcode_type, 16#0D#),
      2674 => to_slv(opcode_type, 16#0B#),
      2675 => to_slv(opcode_type, 16#05#),
      2676 => to_slv(opcode_type, 16#0E#),
      2677 => to_slv(opcode_type, 16#07#),
      2678 => to_slv(opcode_type, 16#09#),
      2679 => to_slv(opcode_type, 16#11#),
      2680 => to_slv(opcode_type, 16#0F#),
      2681 => to_slv(opcode_type, 16#08#),
      2682 => to_slv(opcode_type, 16#0C#),
      2683 => to_slv(opcode_type, 16#10#),
      2684 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#08#),
      2689 => to_slv(opcode_type, 16#07#),
      2690 => to_slv(opcode_type, 16#09#),
      2691 => to_slv(opcode_type, 16#08#),
      2692 => to_slv(opcode_type, 16#C6#),
      2693 => to_slv(opcode_type, 16#0A#),
      2694 => to_slv(opcode_type, 16#08#),
      2695 => to_slv(opcode_type, 16#C5#),
      2696 => to_slv(opcode_type, 16#0E#),
      2697 => to_slv(opcode_type, 16#03#),
      2698 => to_slv(opcode_type, 16#07#),
      2699 => to_slv(opcode_type, 16#10#),
      2700 => to_slv(opcode_type, 16#0D#),
      2701 => to_slv(opcode_type, 16#06#),
      2702 => to_slv(opcode_type, 16#09#),
      2703 => to_slv(opcode_type, 16#09#),
      2704 => to_slv(opcode_type, 16#0E#),
      2705 => to_slv(opcode_type, 16#0C#),
      2706 => to_slv(opcode_type, 16#09#),
      2707 => to_slv(opcode_type, 16#0D#),
      2708 => to_slv(opcode_type, 16#11#),
      2709 => to_slv(opcode_type, 16#06#),
      2710 => to_slv(opcode_type, 16#09#),
      2711 => to_slv(opcode_type, 16#0C#),
      2712 => to_slv(opcode_type, 16#7D#),
      2713 => to_slv(opcode_type, 16#06#),
      2714 => to_slv(opcode_type, 16#A1#),
      2715 => to_slv(opcode_type, 16#0E#),
      2716 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#07#),
      2721 => to_slv(opcode_type, 16#09#),
      2722 => to_slv(opcode_type, 16#03#),
      2723 => to_slv(opcode_type, 16#09#),
      2724 => to_slv(opcode_type, 16#11#),
      2725 => to_slv(opcode_type, 16#0B#),
      2726 => to_slv(opcode_type, 16#06#),
      2727 => to_slv(opcode_type, 16#08#),
      2728 => to_slv(opcode_type, 16#10#),
      2729 => to_slv(opcode_type, 16#0C#),
      2730 => to_slv(opcode_type, 16#08#),
      2731 => to_slv(opcode_type, 16#0E#),
      2732 => to_slv(opcode_type, 16#0F#),
      2733 => to_slv(opcode_type, 16#07#),
      2734 => to_slv(opcode_type, 16#09#),
      2735 => to_slv(opcode_type, 16#06#),
      2736 => to_slv(opcode_type, 16#10#),
      2737 => to_slv(opcode_type, 16#0D#),
      2738 => to_slv(opcode_type, 16#08#),
      2739 => to_slv(opcode_type, 16#0E#),
      2740 => to_slv(opcode_type, 16#0D#),
      2741 => to_slv(opcode_type, 16#06#),
      2742 => to_slv(opcode_type, 16#06#),
      2743 => to_slv(opcode_type, 16#0A#),
      2744 => to_slv(opcode_type, 16#0D#),
      2745 => to_slv(opcode_type, 16#08#),
      2746 => to_slv(opcode_type, 16#7A#),
      2747 => to_slv(opcode_type, 16#10#),
      2748 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#08#),
      2753 => to_slv(opcode_type, 16#07#),
      2754 => to_slv(opcode_type, 16#08#),
      2755 => to_slv(opcode_type, 16#08#),
      2756 => to_slv(opcode_type, 16#11#),
      2757 => to_slv(opcode_type, 16#0F#),
      2758 => to_slv(opcode_type, 16#03#),
      2759 => to_slv(opcode_type, 16#0B#),
      2760 => to_slv(opcode_type, 16#09#),
      2761 => to_slv(opcode_type, 16#02#),
      2762 => to_slv(opcode_type, 16#0C#),
      2763 => to_slv(opcode_type, 16#03#),
      2764 => to_slv(opcode_type, 16#11#),
      2765 => to_slv(opcode_type, 16#07#),
      2766 => to_slv(opcode_type, 16#06#),
      2767 => to_slv(opcode_type, 16#09#),
      2768 => to_slv(opcode_type, 16#0E#),
      2769 => to_slv(opcode_type, 16#0E#),
      2770 => to_slv(opcode_type, 16#07#),
      2771 => to_slv(opcode_type, 16#0A#),
      2772 => to_slv(opcode_type, 16#11#),
      2773 => to_slv(opcode_type, 16#07#),
      2774 => to_slv(opcode_type, 16#07#),
      2775 => to_slv(opcode_type, 16#0C#),
      2776 => to_slv(opcode_type, 16#0E#),
      2777 => to_slv(opcode_type, 16#09#),
      2778 => to_slv(opcode_type, 16#11#),
      2779 => to_slv(opcode_type, 16#0F#),
      2780 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#09#),
      2785 => to_slv(opcode_type, 16#08#),
      2786 => to_slv(opcode_type, 16#02#),
      2787 => to_slv(opcode_type, 16#06#),
      2788 => to_slv(opcode_type, 16#0A#),
      2789 => to_slv(opcode_type, 16#0E#),
      2790 => to_slv(opcode_type, 16#06#),
      2791 => to_slv(opcode_type, 16#06#),
      2792 => to_slv(opcode_type, 16#11#),
      2793 => to_slv(opcode_type, 16#0D#),
      2794 => to_slv(opcode_type, 16#08#),
      2795 => to_slv(opcode_type, 16#0C#),
      2796 => to_slv(opcode_type, 16#11#),
      2797 => to_slv(opcode_type, 16#09#),
      2798 => to_slv(opcode_type, 16#09#),
      2799 => to_slv(opcode_type, 16#09#),
      2800 => to_slv(opcode_type, 16#0B#),
      2801 => to_slv(opcode_type, 16#0A#),
      2802 => to_slv(opcode_type, 16#07#),
      2803 => to_slv(opcode_type, 16#0F#),
      2804 => to_slv(opcode_type, 16#0D#),
      2805 => to_slv(opcode_type, 16#09#),
      2806 => to_slv(opcode_type, 16#09#),
      2807 => to_slv(opcode_type, 16#0A#),
      2808 => to_slv(opcode_type, 16#26#),
      2809 => to_slv(opcode_type, 16#09#),
      2810 => to_slv(opcode_type, 16#0A#),
      2811 => to_slv(opcode_type, 16#EA#),
      2812 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#07#),
      2817 => to_slv(opcode_type, 16#09#),
      2818 => to_slv(opcode_type, 16#01#),
      2819 => to_slv(opcode_type, 16#07#),
      2820 => to_slv(opcode_type, 16#28#),
      2821 => to_slv(opcode_type, 16#11#),
      2822 => to_slv(opcode_type, 16#08#),
      2823 => to_slv(opcode_type, 16#09#),
      2824 => to_slv(opcode_type, 16#A1#),
      2825 => to_slv(opcode_type, 16#0F#),
      2826 => to_slv(opcode_type, 16#08#),
      2827 => to_slv(opcode_type, 16#0A#),
      2828 => to_slv(opcode_type, 16#9A#),
      2829 => to_slv(opcode_type, 16#06#),
      2830 => to_slv(opcode_type, 16#08#),
      2831 => to_slv(opcode_type, 16#07#),
      2832 => to_slv(opcode_type, 16#0D#),
      2833 => to_slv(opcode_type, 16#11#),
      2834 => to_slv(opcode_type, 16#08#),
      2835 => to_slv(opcode_type, 16#0D#),
      2836 => to_slv(opcode_type, 16#10#),
      2837 => to_slv(opcode_type, 16#07#),
      2838 => to_slv(opcode_type, 16#09#),
      2839 => to_slv(opcode_type, 16#0E#),
      2840 => to_slv(opcode_type, 16#11#),
      2841 => to_slv(opcode_type, 16#09#),
      2842 => to_slv(opcode_type, 16#0F#),
      2843 => to_slv(opcode_type, 16#10#),
      2844 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#07#),
      2849 => to_slv(opcode_type, 16#09#),
      2850 => to_slv(opcode_type, 16#01#),
      2851 => to_slv(opcode_type, 16#09#),
      2852 => to_slv(opcode_type, 16#6B#),
      2853 => to_slv(opcode_type, 16#69#),
      2854 => to_slv(opcode_type, 16#08#),
      2855 => to_slv(opcode_type, 16#07#),
      2856 => to_slv(opcode_type, 16#10#),
      2857 => to_slv(opcode_type, 16#0E#),
      2858 => to_slv(opcode_type, 16#08#),
      2859 => to_slv(opcode_type, 16#0E#),
      2860 => to_slv(opcode_type, 16#0E#),
      2861 => to_slv(opcode_type, 16#07#),
      2862 => to_slv(opcode_type, 16#06#),
      2863 => to_slv(opcode_type, 16#06#),
      2864 => to_slv(opcode_type, 16#0A#),
      2865 => to_slv(opcode_type, 16#0A#),
      2866 => to_slv(opcode_type, 16#06#),
      2867 => to_slv(opcode_type, 16#0C#),
      2868 => to_slv(opcode_type, 16#0E#),
      2869 => to_slv(opcode_type, 16#07#),
      2870 => to_slv(opcode_type, 16#07#),
      2871 => to_slv(opcode_type, 16#0F#),
      2872 => to_slv(opcode_type, 16#0D#),
      2873 => to_slv(opcode_type, 16#09#),
      2874 => to_slv(opcode_type, 16#81#),
      2875 => to_slv(opcode_type, 16#0F#),
      2876 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#07#),
      2881 => to_slv(opcode_type, 16#06#),
      2882 => to_slv(opcode_type, 16#08#),
      2883 => to_slv(opcode_type, 16#04#),
      2884 => to_slv(opcode_type, 16#0E#),
      2885 => to_slv(opcode_type, 16#06#),
      2886 => to_slv(opcode_type, 16#0C#),
      2887 => to_slv(opcode_type, 16#0C#),
      2888 => to_slv(opcode_type, 16#06#),
      2889 => to_slv(opcode_type, 16#02#),
      2890 => to_slv(opcode_type, 16#10#),
      2891 => to_slv(opcode_type, 16#05#),
      2892 => to_slv(opcode_type, 16#11#),
      2893 => to_slv(opcode_type, 16#08#),
      2894 => to_slv(opcode_type, 16#09#),
      2895 => to_slv(opcode_type, 16#06#),
      2896 => to_slv(opcode_type, 16#0E#),
      2897 => to_slv(opcode_type, 16#10#),
      2898 => to_slv(opcode_type, 16#06#),
      2899 => to_slv(opcode_type, 16#10#),
      2900 => to_slv(opcode_type, 16#11#),
      2901 => to_slv(opcode_type, 16#09#),
      2902 => to_slv(opcode_type, 16#08#),
      2903 => to_slv(opcode_type, 16#0C#),
      2904 => to_slv(opcode_type, 16#0A#),
      2905 => to_slv(opcode_type, 16#08#),
      2906 => to_slv(opcode_type, 16#0B#),
      2907 => to_slv(opcode_type, 16#76#),
      2908 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#06#),
      2913 => to_slv(opcode_type, 16#07#),
      2914 => to_slv(opcode_type, 16#06#),
      2915 => to_slv(opcode_type, 16#06#),
      2916 => to_slv(opcode_type, 16#0B#),
      2917 => to_slv(opcode_type, 16#0D#),
      2918 => to_slv(opcode_type, 16#06#),
      2919 => to_slv(opcode_type, 16#0F#),
      2920 => to_slv(opcode_type, 16#0A#),
      2921 => to_slv(opcode_type, 16#08#),
      2922 => to_slv(opcode_type, 16#06#),
      2923 => to_slv(opcode_type, 16#10#),
      2924 => to_slv(opcode_type, 16#11#),
      2925 => to_slv(opcode_type, 16#09#),
      2926 => to_slv(opcode_type, 16#0B#),
      2927 => to_slv(opcode_type, 16#0E#),
      2928 => to_slv(opcode_type, 16#09#),
      2929 => to_slv(opcode_type, 16#03#),
      2930 => to_slv(opcode_type, 16#06#),
      2931 => to_slv(opcode_type, 16#0B#),
      2932 => to_slv(opcode_type, 16#0C#),
      2933 => to_slv(opcode_type, 16#07#),
      2934 => to_slv(opcode_type, 16#06#),
      2935 => to_slv(opcode_type, 16#11#),
      2936 => to_slv(opcode_type, 16#0E#),
      2937 => to_slv(opcode_type, 16#09#),
      2938 => to_slv(opcode_type, 16#0F#),
      2939 => to_slv(opcode_type, 16#11#),
      2940 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#06#),
      2945 => to_slv(opcode_type, 16#07#),
      2946 => to_slv(opcode_type, 16#03#),
      2947 => to_slv(opcode_type, 16#09#),
      2948 => to_slv(opcode_type, 16#11#),
      2949 => to_slv(opcode_type, 16#0D#),
      2950 => to_slv(opcode_type, 16#07#),
      2951 => to_slv(opcode_type, 16#07#),
      2952 => to_slv(opcode_type, 16#0E#),
      2953 => to_slv(opcode_type, 16#0C#),
      2954 => to_slv(opcode_type, 16#09#),
      2955 => to_slv(opcode_type, 16#0F#),
      2956 => to_slv(opcode_type, 16#0B#),
      2957 => to_slv(opcode_type, 16#08#),
      2958 => to_slv(opcode_type, 16#08#),
      2959 => to_slv(opcode_type, 16#06#),
      2960 => to_slv(opcode_type, 16#11#),
      2961 => to_slv(opcode_type, 16#0D#),
      2962 => to_slv(opcode_type, 16#09#),
      2963 => to_slv(opcode_type, 16#10#),
      2964 => to_slv(opcode_type, 16#0B#),
      2965 => to_slv(opcode_type, 16#06#),
      2966 => to_slv(opcode_type, 16#06#),
      2967 => to_slv(opcode_type, 16#0F#),
      2968 => to_slv(opcode_type, 16#0B#),
      2969 => to_slv(opcode_type, 16#06#),
      2970 => to_slv(opcode_type, 16#72#),
      2971 => to_slv(opcode_type, 16#0D#),
      2972 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#08#),
      2977 => to_slv(opcode_type, 16#06#),
      2978 => to_slv(opcode_type, 16#04#),
      2979 => to_slv(opcode_type, 16#07#),
      2980 => to_slv(opcode_type, 16#F6#),
      2981 => to_slv(opcode_type, 16#0C#),
      2982 => to_slv(opcode_type, 16#06#),
      2983 => to_slv(opcode_type, 16#08#),
      2984 => to_slv(opcode_type, 16#0F#),
      2985 => to_slv(opcode_type, 16#0A#),
      2986 => to_slv(opcode_type, 16#06#),
      2987 => to_slv(opcode_type, 16#10#),
      2988 => to_slv(opcode_type, 16#72#),
      2989 => to_slv(opcode_type, 16#09#),
      2990 => to_slv(opcode_type, 16#08#),
      2991 => to_slv(opcode_type, 16#06#),
      2992 => to_slv(opcode_type, 16#0D#),
      2993 => to_slv(opcode_type, 16#0C#),
      2994 => to_slv(opcode_type, 16#08#),
      2995 => to_slv(opcode_type, 16#10#),
      2996 => to_slv(opcode_type, 16#0D#),
      2997 => to_slv(opcode_type, 16#09#),
      2998 => to_slv(opcode_type, 16#09#),
      2999 => to_slv(opcode_type, 16#0B#),
      3000 => to_slv(opcode_type, 16#0B#),
      3001 => to_slv(opcode_type, 16#09#),
      3002 => to_slv(opcode_type, 16#0C#),
      3003 => to_slv(opcode_type, 16#0C#),
      3004 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#08#),
      3009 => to_slv(opcode_type, 16#06#),
      3010 => to_slv(opcode_type, 16#07#),
      3011 => to_slv(opcode_type, 16#09#),
      3012 => to_slv(opcode_type, 16#10#),
      3013 => to_slv(opcode_type, 16#0C#),
      3014 => to_slv(opcode_type, 16#09#),
      3015 => to_slv(opcode_type, 16#0B#),
      3016 => to_slv(opcode_type, 16#0A#),
      3017 => to_slv(opcode_type, 16#02#),
      3018 => to_slv(opcode_type, 16#06#),
      3019 => to_slv(opcode_type, 16#0A#),
      3020 => to_slv(opcode_type, 16#0A#),
      3021 => to_slv(opcode_type, 16#09#),
      3022 => to_slv(opcode_type, 16#09#),
      3023 => to_slv(opcode_type, 16#06#),
      3024 => to_slv(opcode_type, 16#0C#),
      3025 => to_slv(opcode_type, 16#10#),
      3026 => to_slv(opcode_type, 16#06#),
      3027 => to_slv(opcode_type, 16#0E#),
      3028 => to_slv(opcode_type, 16#10#),
      3029 => to_slv(opcode_type, 16#08#),
      3030 => to_slv(opcode_type, 16#07#),
      3031 => to_slv(opcode_type, 16#32#),
      3032 => to_slv(opcode_type, 16#0B#),
      3033 => to_slv(opcode_type, 16#08#),
      3034 => to_slv(opcode_type, 16#0B#),
      3035 => to_slv(opcode_type, 16#0C#),
      3036 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#06#),
      3041 => to_slv(opcode_type, 16#08#),
      3042 => to_slv(opcode_type, 16#03#),
      3043 => to_slv(opcode_type, 16#07#),
      3044 => to_slv(opcode_type, 16#0C#),
      3045 => to_slv(opcode_type, 16#0F#),
      3046 => to_slv(opcode_type, 16#08#),
      3047 => to_slv(opcode_type, 16#08#),
      3048 => to_slv(opcode_type, 16#0F#),
      3049 => to_slv(opcode_type, 16#0B#),
      3050 => to_slv(opcode_type, 16#07#),
      3051 => to_slv(opcode_type, 16#0F#),
      3052 => to_slv(opcode_type, 16#0A#),
      3053 => to_slv(opcode_type, 16#09#),
      3054 => to_slv(opcode_type, 16#06#),
      3055 => to_slv(opcode_type, 16#08#),
      3056 => to_slv(opcode_type, 16#0B#),
      3057 => to_slv(opcode_type, 16#0D#),
      3058 => to_slv(opcode_type, 16#09#),
      3059 => to_slv(opcode_type, 16#0B#),
      3060 => to_slv(opcode_type, 16#0E#),
      3061 => to_slv(opcode_type, 16#06#),
      3062 => to_slv(opcode_type, 16#07#),
      3063 => to_slv(opcode_type, 16#0E#),
      3064 => to_slv(opcode_type, 16#0A#),
      3065 => to_slv(opcode_type, 16#08#),
      3066 => to_slv(opcode_type, 16#11#),
      3067 => to_slv(opcode_type, 16#0D#),
      3068 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#08#),
      3073 => to_slv(opcode_type, 16#08#),
      3074 => to_slv(opcode_type, 16#02#),
      3075 => to_slv(opcode_type, 16#07#),
      3076 => to_slv(opcode_type, 16#0B#),
      3077 => to_slv(opcode_type, 16#0C#),
      3078 => to_slv(opcode_type, 16#09#),
      3079 => to_slv(opcode_type, 16#06#),
      3080 => to_slv(opcode_type, 16#0D#),
      3081 => to_slv(opcode_type, 16#0B#),
      3082 => to_slv(opcode_type, 16#09#),
      3083 => to_slv(opcode_type, 16#0D#),
      3084 => to_slv(opcode_type, 16#0B#),
      3085 => to_slv(opcode_type, 16#09#),
      3086 => to_slv(opcode_type, 16#08#),
      3087 => to_slv(opcode_type, 16#06#),
      3088 => to_slv(opcode_type, 16#0C#),
      3089 => to_slv(opcode_type, 16#0A#),
      3090 => to_slv(opcode_type, 16#06#),
      3091 => to_slv(opcode_type, 16#0E#),
      3092 => to_slv(opcode_type, 16#0B#),
      3093 => to_slv(opcode_type, 16#06#),
      3094 => to_slv(opcode_type, 16#09#),
      3095 => to_slv(opcode_type, 16#10#),
      3096 => to_slv(opcode_type, 16#0C#),
      3097 => to_slv(opcode_type, 16#07#),
      3098 => to_slv(opcode_type, 16#0E#),
      3099 => to_slv(opcode_type, 16#0F#),
      3100 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#06#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#04#),
      3107 => to_slv(opcode_type, 16#09#),
      3108 => to_slv(opcode_type, 16#0C#),
      3109 => to_slv(opcode_type, 16#11#),
      3110 => to_slv(opcode_type, 16#08#),
      3111 => to_slv(opcode_type, 16#07#),
      3112 => to_slv(opcode_type, 16#0B#),
      3113 => to_slv(opcode_type, 16#0F#),
      3114 => to_slv(opcode_type, 16#08#),
      3115 => to_slv(opcode_type, 16#0C#),
      3116 => to_slv(opcode_type, 16#0A#),
      3117 => to_slv(opcode_type, 16#09#),
      3118 => to_slv(opcode_type, 16#06#),
      3119 => to_slv(opcode_type, 16#06#),
      3120 => to_slv(opcode_type, 16#10#),
      3121 => to_slv(opcode_type, 16#0A#),
      3122 => to_slv(opcode_type, 16#07#),
      3123 => to_slv(opcode_type, 16#10#),
      3124 => to_slv(opcode_type, 16#0C#),
      3125 => to_slv(opcode_type, 16#09#),
      3126 => to_slv(opcode_type, 16#06#),
      3127 => to_slv(opcode_type, 16#0C#),
      3128 => to_slv(opcode_type, 16#0D#),
      3129 => to_slv(opcode_type, 16#08#),
      3130 => to_slv(opcode_type, 16#12#),
      3131 => to_slv(opcode_type, 16#0C#),
      3132 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#09#),
      3137 => to_slv(opcode_type, 16#09#),
      3138 => to_slv(opcode_type, 16#09#),
      3139 => to_slv(opcode_type, 16#09#),
      3140 => to_slv(opcode_type, 16#0A#),
      3141 => to_slv(opcode_type, 16#B0#),
      3142 => to_slv(opcode_type, 16#05#),
      3143 => to_slv(opcode_type, 16#10#),
      3144 => to_slv(opcode_type, 16#07#),
      3145 => to_slv(opcode_type, 16#09#),
      3146 => to_slv(opcode_type, 16#0D#),
      3147 => to_slv(opcode_type, 16#0B#),
      3148 => to_slv(opcode_type, 16#04#),
      3149 => to_slv(opcode_type, 16#0C#),
      3150 => to_slv(opcode_type, 16#09#),
      3151 => to_slv(opcode_type, 16#06#),
      3152 => to_slv(opcode_type, 16#06#),
      3153 => to_slv(opcode_type, 16#0F#),
      3154 => to_slv(opcode_type, 16#11#),
      3155 => to_slv(opcode_type, 16#09#),
      3156 => to_slv(opcode_type, 16#10#),
      3157 => to_slv(opcode_type, 16#10#),
      3158 => to_slv(opcode_type, 16#09#),
      3159 => to_slv(opcode_type, 16#02#),
      3160 => to_slv(opcode_type, 16#0B#),
      3161 => to_slv(opcode_type, 16#06#),
      3162 => to_slv(opcode_type, 16#0C#),
      3163 => to_slv(opcode_type, 16#0A#),
      3164 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#08#),
      3169 => to_slv(opcode_type, 16#07#),
      3170 => to_slv(opcode_type, 16#07#),
      3171 => to_slv(opcode_type, 16#06#),
      3172 => to_slv(opcode_type, 16#10#),
      3173 => to_slv(opcode_type, 16#0D#),
      3174 => to_slv(opcode_type, 16#04#),
      3175 => to_slv(opcode_type, 16#0F#),
      3176 => to_slv(opcode_type, 16#06#),
      3177 => to_slv(opcode_type, 16#01#),
      3178 => to_slv(opcode_type, 16#0E#),
      3179 => to_slv(opcode_type, 16#08#),
      3180 => to_slv(opcode_type, 16#0D#),
      3181 => to_slv(opcode_type, 16#0E#),
      3182 => to_slv(opcode_type, 16#08#),
      3183 => to_slv(opcode_type, 16#07#),
      3184 => to_slv(opcode_type, 16#05#),
      3185 => to_slv(opcode_type, 16#0E#),
      3186 => to_slv(opcode_type, 16#07#),
      3187 => to_slv(opcode_type, 16#11#),
      3188 => to_slv(opcode_type, 16#11#),
      3189 => to_slv(opcode_type, 16#09#),
      3190 => to_slv(opcode_type, 16#09#),
      3191 => to_slv(opcode_type, 16#0E#),
      3192 => to_slv(opcode_type, 16#0F#),
      3193 => to_slv(opcode_type, 16#09#),
      3194 => to_slv(opcode_type, 16#0D#),
      3195 => to_slv(opcode_type, 16#0C#),
      3196 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#08#),
      3201 => to_slv(opcode_type, 16#07#),
      3202 => to_slv(opcode_type, 16#03#),
      3203 => to_slv(opcode_type, 16#07#),
      3204 => to_slv(opcode_type, 16#0F#),
      3205 => to_slv(opcode_type, 16#10#),
      3206 => to_slv(opcode_type, 16#07#),
      3207 => to_slv(opcode_type, 16#08#),
      3208 => to_slv(opcode_type, 16#0E#),
      3209 => to_slv(opcode_type, 16#93#),
      3210 => to_slv(opcode_type, 16#08#),
      3211 => to_slv(opcode_type, 16#11#),
      3212 => to_slv(opcode_type, 16#0E#),
      3213 => to_slv(opcode_type, 16#07#),
      3214 => to_slv(opcode_type, 16#08#),
      3215 => to_slv(opcode_type, 16#09#),
      3216 => to_slv(opcode_type, 16#0D#),
      3217 => to_slv(opcode_type, 16#10#),
      3218 => to_slv(opcode_type, 16#08#),
      3219 => to_slv(opcode_type, 16#0C#),
      3220 => to_slv(opcode_type, 16#0A#),
      3221 => to_slv(opcode_type, 16#07#),
      3222 => to_slv(opcode_type, 16#06#),
      3223 => to_slv(opcode_type, 16#0C#),
      3224 => to_slv(opcode_type, 16#0E#),
      3225 => to_slv(opcode_type, 16#08#),
      3226 => to_slv(opcode_type, 16#11#),
      3227 => to_slv(opcode_type, 16#8B#),
      3228 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#07#),
      3233 => to_slv(opcode_type, 16#08#),
      3234 => to_slv(opcode_type, 16#04#),
      3235 => to_slv(opcode_type, 16#08#),
      3236 => to_slv(opcode_type, 16#0A#),
      3237 => to_slv(opcode_type, 16#11#),
      3238 => to_slv(opcode_type, 16#08#),
      3239 => to_slv(opcode_type, 16#07#),
      3240 => to_slv(opcode_type, 16#A5#),
      3241 => to_slv(opcode_type, 16#A9#),
      3242 => to_slv(opcode_type, 16#06#),
      3243 => to_slv(opcode_type, 16#0D#),
      3244 => to_slv(opcode_type, 16#0F#),
      3245 => to_slv(opcode_type, 16#07#),
      3246 => to_slv(opcode_type, 16#06#),
      3247 => to_slv(opcode_type, 16#09#),
      3248 => to_slv(opcode_type, 16#0E#),
      3249 => to_slv(opcode_type, 16#0B#),
      3250 => to_slv(opcode_type, 16#08#),
      3251 => to_slv(opcode_type, 16#0A#),
      3252 => to_slv(opcode_type, 16#0C#),
      3253 => to_slv(opcode_type, 16#08#),
      3254 => to_slv(opcode_type, 16#08#),
      3255 => to_slv(opcode_type, 16#0B#),
      3256 => to_slv(opcode_type, 16#0E#),
      3257 => to_slv(opcode_type, 16#08#),
      3258 => to_slv(opcode_type, 16#0D#),
      3259 => to_slv(opcode_type, 16#0E#),
      3260 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#06#),
      3265 => to_slv(opcode_type, 16#06#),
      3266 => to_slv(opcode_type, 16#05#),
      3267 => to_slv(opcode_type, 16#08#),
      3268 => to_slv(opcode_type, 16#0A#),
      3269 => to_slv(opcode_type, 16#0B#),
      3270 => to_slv(opcode_type, 16#06#),
      3271 => to_slv(opcode_type, 16#09#),
      3272 => to_slv(opcode_type, 16#0C#),
      3273 => to_slv(opcode_type, 16#0B#),
      3274 => to_slv(opcode_type, 16#09#),
      3275 => to_slv(opcode_type, 16#11#),
      3276 => to_slv(opcode_type, 16#0A#),
      3277 => to_slv(opcode_type, 16#07#),
      3278 => to_slv(opcode_type, 16#08#),
      3279 => to_slv(opcode_type, 16#09#),
      3280 => to_slv(opcode_type, 16#0D#),
      3281 => to_slv(opcode_type, 16#0A#),
      3282 => to_slv(opcode_type, 16#09#),
      3283 => to_slv(opcode_type, 16#0A#),
      3284 => to_slv(opcode_type, 16#0F#),
      3285 => to_slv(opcode_type, 16#09#),
      3286 => to_slv(opcode_type, 16#07#),
      3287 => to_slv(opcode_type, 16#11#),
      3288 => to_slv(opcode_type, 16#11#),
      3289 => to_slv(opcode_type, 16#06#),
      3290 => to_slv(opcode_type, 16#1A#),
      3291 => to_slv(opcode_type, 16#0E#),
      3292 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#07#),
      3297 => to_slv(opcode_type, 16#07#),
      3298 => to_slv(opcode_type, 16#02#),
      3299 => to_slv(opcode_type, 16#08#),
      3300 => to_slv(opcode_type, 16#0E#),
      3301 => to_slv(opcode_type, 16#11#),
      3302 => to_slv(opcode_type, 16#08#),
      3303 => to_slv(opcode_type, 16#06#),
      3304 => to_slv(opcode_type, 16#0C#),
      3305 => to_slv(opcode_type, 16#0F#),
      3306 => to_slv(opcode_type, 16#09#),
      3307 => to_slv(opcode_type, 16#0B#),
      3308 => to_slv(opcode_type, 16#0E#),
      3309 => to_slv(opcode_type, 16#09#),
      3310 => to_slv(opcode_type, 16#09#),
      3311 => to_slv(opcode_type, 16#06#),
      3312 => to_slv(opcode_type, 16#0A#),
      3313 => to_slv(opcode_type, 16#0C#),
      3314 => to_slv(opcode_type, 16#06#),
      3315 => to_slv(opcode_type, 16#0D#),
      3316 => to_slv(opcode_type, 16#10#),
      3317 => to_slv(opcode_type, 16#09#),
      3318 => to_slv(opcode_type, 16#08#),
      3319 => to_slv(opcode_type, 16#0B#),
      3320 => to_slv(opcode_type, 16#0D#),
      3321 => to_slv(opcode_type, 16#07#),
      3322 => to_slv(opcode_type, 16#0A#),
      3323 => to_slv(opcode_type, 16#0F#),
      3324 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#07#),
      3329 => to_slv(opcode_type, 16#07#),
      3330 => to_slv(opcode_type, 16#08#),
      3331 => to_slv(opcode_type, 16#02#),
      3332 => to_slv(opcode_type, 16#0E#),
      3333 => to_slv(opcode_type, 16#03#),
      3334 => to_slv(opcode_type, 16#0C#),
      3335 => to_slv(opcode_type, 16#06#),
      3336 => to_slv(opcode_type, 16#08#),
      3337 => to_slv(opcode_type, 16#0B#),
      3338 => to_slv(opcode_type, 16#0A#),
      3339 => to_slv(opcode_type, 16#09#),
      3340 => to_slv(opcode_type, 16#69#),
      3341 => to_slv(opcode_type, 16#10#),
      3342 => to_slv(opcode_type, 16#06#),
      3343 => to_slv(opcode_type, 16#06#),
      3344 => to_slv(opcode_type, 16#04#),
      3345 => to_slv(opcode_type, 16#D0#),
      3346 => to_slv(opcode_type, 16#09#),
      3347 => to_slv(opcode_type, 16#0F#),
      3348 => to_slv(opcode_type, 16#0A#),
      3349 => to_slv(opcode_type, 16#08#),
      3350 => to_slv(opcode_type, 16#07#),
      3351 => to_slv(opcode_type, 16#0B#),
      3352 => to_slv(opcode_type, 16#0E#),
      3353 => to_slv(opcode_type, 16#09#),
      3354 => to_slv(opcode_type, 16#0A#),
      3355 => to_slv(opcode_type, 16#0F#),
      3356 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#08#),
      3361 => to_slv(opcode_type, 16#07#),
      3362 => to_slv(opcode_type, 16#05#),
      3363 => to_slv(opcode_type, 16#06#),
      3364 => to_slv(opcode_type, 16#0F#),
      3365 => to_slv(opcode_type, 16#0E#),
      3366 => to_slv(opcode_type, 16#06#),
      3367 => to_slv(opcode_type, 16#06#),
      3368 => to_slv(opcode_type, 16#EF#),
      3369 => to_slv(opcode_type, 16#10#),
      3370 => to_slv(opcode_type, 16#07#),
      3371 => to_slv(opcode_type, 16#10#),
      3372 => to_slv(opcode_type, 16#0A#),
      3373 => to_slv(opcode_type, 16#06#),
      3374 => to_slv(opcode_type, 16#09#),
      3375 => to_slv(opcode_type, 16#08#),
      3376 => to_slv(opcode_type, 16#0E#),
      3377 => to_slv(opcode_type, 16#0C#),
      3378 => to_slv(opcode_type, 16#08#),
      3379 => to_slv(opcode_type, 16#0F#),
      3380 => to_slv(opcode_type, 16#0A#),
      3381 => to_slv(opcode_type, 16#07#),
      3382 => to_slv(opcode_type, 16#09#),
      3383 => to_slv(opcode_type, 16#11#),
      3384 => to_slv(opcode_type, 16#0D#),
      3385 => to_slv(opcode_type, 16#07#),
      3386 => to_slv(opcode_type, 16#0F#),
      3387 => to_slv(opcode_type, 16#0B#),
      3388 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#08#),
      3393 => to_slv(opcode_type, 16#08#),
      3394 => to_slv(opcode_type, 16#05#),
      3395 => to_slv(opcode_type, 16#06#),
      3396 => to_slv(opcode_type, 16#0B#),
      3397 => to_slv(opcode_type, 16#12#),
      3398 => to_slv(opcode_type, 16#06#),
      3399 => to_slv(opcode_type, 16#07#),
      3400 => to_slv(opcode_type, 16#0E#),
      3401 => to_slv(opcode_type, 16#0C#),
      3402 => to_slv(opcode_type, 16#09#),
      3403 => to_slv(opcode_type, 16#11#),
      3404 => to_slv(opcode_type, 16#11#),
      3405 => to_slv(opcode_type, 16#08#),
      3406 => to_slv(opcode_type, 16#08#),
      3407 => to_slv(opcode_type, 16#09#),
      3408 => to_slv(opcode_type, 16#0B#),
      3409 => to_slv(opcode_type, 16#11#),
      3410 => to_slv(opcode_type, 16#06#),
      3411 => to_slv(opcode_type, 16#11#),
      3412 => to_slv(opcode_type, 16#0A#),
      3413 => to_slv(opcode_type, 16#09#),
      3414 => to_slv(opcode_type, 16#06#),
      3415 => to_slv(opcode_type, 16#11#),
      3416 => to_slv(opcode_type, 16#61#),
      3417 => to_slv(opcode_type, 16#08#),
      3418 => to_slv(opcode_type, 16#0D#),
      3419 => to_slv(opcode_type, 16#E1#),
      3420 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#08#),
      3425 => to_slv(opcode_type, 16#08#),
      3426 => to_slv(opcode_type, 16#04#),
      3427 => to_slv(opcode_type, 16#09#),
      3428 => to_slv(opcode_type, 16#0E#),
      3429 => to_slv(opcode_type, 16#11#),
      3430 => to_slv(opcode_type, 16#07#),
      3431 => to_slv(opcode_type, 16#09#),
      3432 => to_slv(opcode_type, 16#0B#),
      3433 => to_slv(opcode_type, 16#69#),
      3434 => to_slv(opcode_type, 16#07#),
      3435 => to_slv(opcode_type, 16#10#),
      3436 => to_slv(opcode_type, 16#0B#),
      3437 => to_slv(opcode_type, 16#08#),
      3438 => to_slv(opcode_type, 16#08#),
      3439 => to_slv(opcode_type, 16#07#),
      3440 => to_slv(opcode_type, 16#0D#),
      3441 => to_slv(opcode_type, 16#0A#),
      3442 => to_slv(opcode_type, 16#06#),
      3443 => to_slv(opcode_type, 16#0E#),
      3444 => to_slv(opcode_type, 16#0F#),
      3445 => to_slv(opcode_type, 16#08#),
      3446 => to_slv(opcode_type, 16#08#),
      3447 => to_slv(opcode_type, 16#0F#),
      3448 => to_slv(opcode_type, 16#0B#),
      3449 => to_slv(opcode_type, 16#07#),
      3450 => to_slv(opcode_type, 16#0C#),
      3451 => to_slv(opcode_type, 16#0F#),
      3452 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#09#),
      3457 => to_slv(opcode_type, 16#07#),
      3458 => to_slv(opcode_type, 16#04#),
      3459 => to_slv(opcode_type, 16#09#),
      3460 => to_slv(opcode_type, 16#10#),
      3461 => to_slv(opcode_type, 16#0F#),
      3462 => to_slv(opcode_type, 16#07#),
      3463 => to_slv(opcode_type, 16#09#),
      3464 => to_slv(opcode_type, 16#0C#),
      3465 => to_slv(opcode_type, 16#11#),
      3466 => to_slv(opcode_type, 16#09#),
      3467 => to_slv(opcode_type, 16#0E#),
      3468 => to_slv(opcode_type, 16#5E#),
      3469 => to_slv(opcode_type, 16#09#),
      3470 => to_slv(opcode_type, 16#09#),
      3471 => to_slv(opcode_type, 16#09#),
      3472 => to_slv(opcode_type, 16#3F#),
      3473 => to_slv(opcode_type, 16#0E#),
      3474 => to_slv(opcode_type, 16#07#),
      3475 => to_slv(opcode_type, 16#11#),
      3476 => to_slv(opcode_type, 16#11#),
      3477 => to_slv(opcode_type, 16#09#),
      3478 => to_slv(opcode_type, 16#06#),
      3479 => to_slv(opcode_type, 16#11#),
      3480 => to_slv(opcode_type, 16#10#),
      3481 => to_slv(opcode_type, 16#09#),
      3482 => to_slv(opcode_type, 16#0D#),
      3483 => to_slv(opcode_type, 16#0C#),
      3484 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#09#),
      3489 => to_slv(opcode_type, 16#07#),
      3490 => to_slv(opcode_type, 16#06#),
      3491 => to_slv(opcode_type, 16#01#),
      3492 => to_slv(opcode_type, 16#0F#),
      3493 => to_slv(opcode_type, 16#02#),
      3494 => to_slv(opcode_type, 16#17#),
      3495 => to_slv(opcode_type, 16#06#),
      3496 => to_slv(opcode_type, 16#05#),
      3497 => to_slv(opcode_type, 16#0E#),
      3498 => to_slv(opcode_type, 16#06#),
      3499 => to_slv(opcode_type, 16#7B#),
      3500 => to_slv(opcode_type, 16#0D#),
      3501 => to_slv(opcode_type, 16#07#),
      3502 => to_slv(opcode_type, 16#08#),
      3503 => to_slv(opcode_type, 16#08#),
      3504 => to_slv(opcode_type, 16#0D#),
      3505 => to_slv(opcode_type, 16#0A#),
      3506 => to_slv(opcode_type, 16#07#),
      3507 => to_slv(opcode_type, 16#0E#),
      3508 => to_slv(opcode_type, 16#0E#),
      3509 => to_slv(opcode_type, 16#07#),
      3510 => to_slv(opcode_type, 16#06#),
      3511 => to_slv(opcode_type, 16#0F#),
      3512 => to_slv(opcode_type, 16#0B#),
      3513 => to_slv(opcode_type, 16#09#),
      3514 => to_slv(opcode_type, 16#11#),
      3515 => to_slv(opcode_type, 16#11#),
      3516 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#06#),
      3521 => to_slv(opcode_type, 16#06#),
      3522 => to_slv(opcode_type, 16#02#),
      3523 => to_slv(opcode_type, 16#06#),
      3524 => to_slv(opcode_type, 16#0A#),
      3525 => to_slv(opcode_type, 16#0F#),
      3526 => to_slv(opcode_type, 16#08#),
      3527 => to_slv(opcode_type, 16#06#),
      3528 => to_slv(opcode_type, 16#10#),
      3529 => to_slv(opcode_type, 16#0E#),
      3530 => to_slv(opcode_type, 16#07#),
      3531 => to_slv(opcode_type, 16#0A#),
      3532 => to_slv(opcode_type, 16#0A#),
      3533 => to_slv(opcode_type, 16#09#),
      3534 => to_slv(opcode_type, 16#06#),
      3535 => to_slv(opcode_type, 16#09#),
      3536 => to_slv(opcode_type, 16#10#),
      3537 => to_slv(opcode_type, 16#0C#),
      3538 => to_slv(opcode_type, 16#06#),
      3539 => to_slv(opcode_type, 16#0D#),
      3540 => to_slv(opcode_type, 16#0E#),
      3541 => to_slv(opcode_type, 16#09#),
      3542 => to_slv(opcode_type, 16#09#),
      3543 => to_slv(opcode_type, 16#11#),
      3544 => to_slv(opcode_type, 16#0D#),
      3545 => to_slv(opcode_type, 16#08#),
      3546 => to_slv(opcode_type, 16#3D#),
      3547 => to_slv(opcode_type, 16#0E#),
      3548 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#06#),
      3553 => to_slv(opcode_type, 16#09#),
      3554 => to_slv(opcode_type, 16#09#),
      3555 => to_slv(opcode_type, 16#07#),
      3556 => to_slv(opcode_type, 16#0C#),
      3557 => to_slv(opcode_type, 16#47#),
      3558 => to_slv(opcode_type, 16#07#),
      3559 => to_slv(opcode_type, 16#0D#),
      3560 => to_slv(opcode_type, 16#11#),
      3561 => to_slv(opcode_type, 16#02#),
      3562 => to_slv(opcode_type, 16#09#),
      3563 => to_slv(opcode_type, 16#0E#),
      3564 => to_slv(opcode_type, 16#C7#),
      3565 => to_slv(opcode_type, 16#08#),
      3566 => to_slv(opcode_type, 16#07#),
      3567 => to_slv(opcode_type, 16#07#),
      3568 => to_slv(opcode_type, 16#10#),
      3569 => to_slv(opcode_type, 16#0D#),
      3570 => to_slv(opcode_type, 16#08#),
      3571 => to_slv(opcode_type, 16#0B#),
      3572 => to_slv(opcode_type, 16#0B#),
      3573 => to_slv(opcode_type, 16#06#),
      3574 => to_slv(opcode_type, 16#07#),
      3575 => to_slv(opcode_type, 16#0D#),
      3576 => to_slv(opcode_type, 16#4C#),
      3577 => to_slv(opcode_type, 16#09#),
      3578 => to_slv(opcode_type, 16#9C#),
      3579 => to_slv(opcode_type, 16#0F#),
      3580 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#06#),
      3585 => to_slv(opcode_type, 16#07#),
      3586 => to_slv(opcode_type, 16#05#),
      3587 => to_slv(opcode_type, 16#09#),
      3588 => to_slv(opcode_type, 16#0D#),
      3589 => to_slv(opcode_type, 16#0A#),
      3590 => to_slv(opcode_type, 16#09#),
      3591 => to_slv(opcode_type, 16#09#),
      3592 => to_slv(opcode_type, 16#6C#),
      3593 => to_slv(opcode_type, 16#0D#),
      3594 => to_slv(opcode_type, 16#07#),
      3595 => to_slv(opcode_type, 16#10#),
      3596 => to_slv(opcode_type, 16#0A#),
      3597 => to_slv(opcode_type, 16#07#),
      3598 => to_slv(opcode_type, 16#07#),
      3599 => to_slv(opcode_type, 16#06#),
      3600 => to_slv(opcode_type, 16#0B#),
      3601 => to_slv(opcode_type, 16#0D#),
      3602 => to_slv(opcode_type, 16#09#),
      3603 => to_slv(opcode_type, 16#A5#),
      3604 => to_slv(opcode_type, 16#0F#),
      3605 => to_slv(opcode_type, 16#08#),
      3606 => to_slv(opcode_type, 16#07#),
      3607 => to_slv(opcode_type, 16#0F#),
      3608 => to_slv(opcode_type, 16#0E#),
      3609 => to_slv(opcode_type, 16#06#),
      3610 => to_slv(opcode_type, 16#0E#),
      3611 => to_slv(opcode_type, 16#11#),
      3612 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#06#),
      3617 => to_slv(opcode_type, 16#07#),
      3618 => to_slv(opcode_type, 16#09#),
      3619 => to_slv(opcode_type, 16#01#),
      3620 => to_slv(opcode_type, 16#0A#),
      3621 => to_slv(opcode_type, 16#09#),
      3622 => to_slv(opcode_type, 16#11#),
      3623 => to_slv(opcode_type, 16#0D#),
      3624 => to_slv(opcode_type, 16#09#),
      3625 => to_slv(opcode_type, 16#07#),
      3626 => to_slv(opcode_type, 16#CC#),
      3627 => to_slv(opcode_type, 16#0E#),
      3628 => to_slv(opcode_type, 16#04#),
      3629 => to_slv(opcode_type, 16#11#),
      3630 => to_slv(opcode_type, 16#07#),
      3631 => to_slv(opcode_type, 16#09#),
      3632 => to_slv(opcode_type, 16#08#),
      3633 => to_slv(opcode_type, 16#11#),
      3634 => to_slv(opcode_type, 16#10#),
      3635 => to_slv(opcode_type, 16#08#),
      3636 => to_slv(opcode_type, 16#0D#),
      3637 => to_slv(opcode_type, 16#0C#),
      3638 => to_slv(opcode_type, 16#08#),
      3639 => to_slv(opcode_type, 16#06#),
      3640 => to_slv(opcode_type, 16#0E#),
      3641 => to_slv(opcode_type, 16#11#),
      3642 => to_slv(opcode_type, 16#02#),
      3643 => to_slv(opcode_type, 16#0D#),
      3644 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#08#),
      3649 => to_slv(opcode_type, 16#09#),
      3650 => to_slv(opcode_type, 16#06#),
      3651 => to_slv(opcode_type, 16#08#),
      3652 => to_slv(opcode_type, 16#10#),
      3653 => to_slv(opcode_type, 16#65#),
      3654 => to_slv(opcode_type, 16#04#),
      3655 => to_slv(opcode_type, 16#0C#),
      3656 => to_slv(opcode_type, 16#09#),
      3657 => to_slv(opcode_type, 16#09#),
      3658 => to_slv(opcode_type, 16#0A#),
      3659 => to_slv(opcode_type, 16#0C#),
      3660 => to_slv(opcode_type, 16#09#),
      3661 => to_slv(opcode_type, 16#0E#),
      3662 => to_slv(opcode_type, 16#0E#),
      3663 => to_slv(opcode_type, 16#07#),
      3664 => to_slv(opcode_type, 16#08#),
      3665 => to_slv(opcode_type, 16#04#),
      3666 => to_slv(opcode_type, 16#11#),
      3667 => to_slv(opcode_type, 16#09#),
      3668 => to_slv(opcode_type, 16#11#),
      3669 => to_slv(opcode_type, 16#0C#),
      3670 => to_slv(opcode_type, 16#07#),
      3671 => to_slv(opcode_type, 16#08#),
      3672 => to_slv(opcode_type, 16#11#),
      3673 => to_slv(opcode_type, 16#0E#),
      3674 => to_slv(opcode_type, 16#05#),
      3675 => to_slv(opcode_type, 16#0E#),
      3676 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#06#),
      3681 => to_slv(opcode_type, 16#08#),
      3682 => to_slv(opcode_type, 16#04#),
      3683 => to_slv(opcode_type, 16#08#),
      3684 => to_slv(opcode_type, 16#0C#),
      3685 => to_slv(opcode_type, 16#0D#),
      3686 => to_slv(opcode_type, 16#09#),
      3687 => to_slv(opcode_type, 16#09#),
      3688 => to_slv(opcode_type, 16#F4#),
      3689 => to_slv(opcode_type, 16#0C#),
      3690 => to_slv(opcode_type, 16#09#),
      3691 => to_slv(opcode_type, 16#0B#),
      3692 => to_slv(opcode_type, 16#0E#),
      3693 => to_slv(opcode_type, 16#08#),
      3694 => to_slv(opcode_type, 16#08#),
      3695 => to_slv(opcode_type, 16#06#),
      3696 => to_slv(opcode_type, 16#10#),
      3697 => to_slv(opcode_type, 16#B6#),
      3698 => to_slv(opcode_type, 16#06#),
      3699 => to_slv(opcode_type, 16#0E#),
      3700 => to_slv(opcode_type, 16#0C#),
      3701 => to_slv(opcode_type, 16#09#),
      3702 => to_slv(opcode_type, 16#09#),
      3703 => to_slv(opcode_type, 16#11#),
      3704 => to_slv(opcode_type, 16#11#),
      3705 => to_slv(opcode_type, 16#07#),
      3706 => to_slv(opcode_type, 16#0C#),
      3707 => to_slv(opcode_type, 16#0D#),
      3708 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#09#),
      3713 => to_slv(opcode_type, 16#07#),
      3714 => to_slv(opcode_type, 16#09#),
      3715 => to_slv(opcode_type, 16#07#),
      3716 => to_slv(opcode_type, 16#0B#),
      3717 => to_slv(opcode_type, 16#0A#),
      3718 => to_slv(opcode_type, 16#09#),
      3719 => to_slv(opcode_type, 16#10#),
      3720 => to_slv(opcode_type, 16#10#),
      3721 => to_slv(opcode_type, 16#09#),
      3722 => to_slv(opcode_type, 16#07#),
      3723 => to_slv(opcode_type, 16#10#),
      3724 => to_slv(opcode_type, 16#0A#),
      3725 => to_slv(opcode_type, 16#09#),
      3726 => to_slv(opcode_type, 16#0D#),
      3727 => to_slv(opcode_type, 16#0D#),
      3728 => to_slv(opcode_type, 16#07#),
      3729 => to_slv(opcode_type, 16#03#),
      3730 => to_slv(opcode_type, 16#08#),
      3731 => to_slv(opcode_type, 16#0B#),
      3732 => to_slv(opcode_type, 16#0A#),
      3733 => to_slv(opcode_type, 16#08#),
      3734 => to_slv(opcode_type, 16#07#),
      3735 => to_slv(opcode_type, 16#0C#),
      3736 => to_slv(opcode_type, 16#0A#),
      3737 => to_slv(opcode_type, 16#06#),
      3738 => to_slv(opcode_type, 16#0E#),
      3739 => to_slv(opcode_type, 16#AB#),
      3740 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#06#),
      3745 => to_slv(opcode_type, 16#08#),
      3746 => to_slv(opcode_type, 16#03#),
      3747 => to_slv(opcode_type, 16#08#),
      3748 => to_slv(opcode_type, 16#0A#),
      3749 => to_slv(opcode_type, 16#0D#),
      3750 => to_slv(opcode_type, 16#07#),
      3751 => to_slv(opcode_type, 16#07#),
      3752 => to_slv(opcode_type, 16#39#),
      3753 => to_slv(opcode_type, 16#11#),
      3754 => to_slv(opcode_type, 16#07#),
      3755 => to_slv(opcode_type, 16#0E#),
      3756 => to_slv(opcode_type, 16#24#),
      3757 => to_slv(opcode_type, 16#08#),
      3758 => to_slv(opcode_type, 16#09#),
      3759 => to_slv(opcode_type, 16#08#),
      3760 => to_slv(opcode_type, 16#10#),
      3761 => to_slv(opcode_type, 16#10#),
      3762 => to_slv(opcode_type, 16#09#),
      3763 => to_slv(opcode_type, 16#0B#),
      3764 => to_slv(opcode_type, 16#0D#),
      3765 => to_slv(opcode_type, 16#09#),
      3766 => to_slv(opcode_type, 16#07#),
      3767 => to_slv(opcode_type, 16#0A#),
      3768 => to_slv(opcode_type, 16#0E#),
      3769 => to_slv(opcode_type, 16#06#),
      3770 => to_slv(opcode_type, 16#0D#),
      3771 => to_slv(opcode_type, 16#0D#),
      3772 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#06#),
      3777 => to_slv(opcode_type, 16#08#),
      3778 => to_slv(opcode_type, 16#01#),
      3779 => to_slv(opcode_type, 16#07#),
      3780 => to_slv(opcode_type, 16#89#),
      3781 => to_slv(opcode_type, 16#10#),
      3782 => to_slv(opcode_type, 16#08#),
      3783 => to_slv(opcode_type, 16#06#),
      3784 => to_slv(opcode_type, 16#0F#),
      3785 => to_slv(opcode_type, 16#11#),
      3786 => to_slv(opcode_type, 16#08#),
      3787 => to_slv(opcode_type, 16#0A#),
      3788 => to_slv(opcode_type, 16#11#),
      3789 => to_slv(opcode_type, 16#07#),
      3790 => to_slv(opcode_type, 16#08#),
      3791 => to_slv(opcode_type, 16#06#),
      3792 => to_slv(opcode_type, 16#0D#),
      3793 => to_slv(opcode_type, 16#0E#),
      3794 => to_slv(opcode_type, 16#09#),
      3795 => to_slv(opcode_type, 16#0E#),
      3796 => to_slv(opcode_type, 16#F5#),
      3797 => to_slv(opcode_type, 16#09#),
      3798 => to_slv(opcode_type, 16#09#),
      3799 => to_slv(opcode_type, 16#F0#),
      3800 => to_slv(opcode_type, 16#0D#),
      3801 => to_slv(opcode_type, 16#09#),
      3802 => to_slv(opcode_type, 16#0E#),
      3803 => to_slv(opcode_type, 16#11#),
      3804 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#09#),
      3809 => to_slv(opcode_type, 16#08#),
      3810 => to_slv(opcode_type, 16#05#),
      3811 => to_slv(opcode_type, 16#08#),
      3812 => to_slv(opcode_type, 16#0E#),
      3813 => to_slv(opcode_type, 16#10#),
      3814 => to_slv(opcode_type, 16#08#),
      3815 => to_slv(opcode_type, 16#08#),
      3816 => to_slv(opcode_type, 16#0B#),
      3817 => to_slv(opcode_type, 16#0D#),
      3818 => to_slv(opcode_type, 16#08#),
      3819 => to_slv(opcode_type, 16#0E#),
      3820 => to_slv(opcode_type, 16#0B#),
      3821 => to_slv(opcode_type, 16#06#),
      3822 => to_slv(opcode_type, 16#08#),
      3823 => to_slv(opcode_type, 16#06#),
      3824 => to_slv(opcode_type, 16#0E#),
      3825 => to_slv(opcode_type, 16#0C#),
      3826 => to_slv(opcode_type, 16#08#),
      3827 => to_slv(opcode_type, 16#0F#),
      3828 => to_slv(opcode_type, 16#0D#),
      3829 => to_slv(opcode_type, 16#09#),
      3830 => to_slv(opcode_type, 16#09#),
      3831 => to_slv(opcode_type, 16#0C#),
      3832 => to_slv(opcode_type, 16#0F#),
      3833 => to_slv(opcode_type, 16#08#),
      3834 => to_slv(opcode_type, 16#CD#),
      3835 => to_slv(opcode_type, 16#11#),
      3836 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#06#),
      3841 => to_slv(opcode_type, 16#09#),
      3842 => to_slv(opcode_type, 16#05#),
      3843 => to_slv(opcode_type, 16#06#),
      3844 => to_slv(opcode_type, 16#0F#),
      3845 => to_slv(opcode_type, 16#10#),
      3846 => to_slv(opcode_type, 16#09#),
      3847 => to_slv(opcode_type, 16#07#),
      3848 => to_slv(opcode_type, 16#11#),
      3849 => to_slv(opcode_type, 16#FE#),
      3850 => to_slv(opcode_type, 16#06#),
      3851 => to_slv(opcode_type, 16#0F#),
      3852 => to_slv(opcode_type, 16#0A#),
      3853 => to_slv(opcode_type, 16#09#),
      3854 => to_slv(opcode_type, 16#07#),
      3855 => to_slv(opcode_type, 16#09#),
      3856 => to_slv(opcode_type, 16#10#),
      3857 => to_slv(opcode_type, 16#0E#),
      3858 => to_slv(opcode_type, 16#06#),
      3859 => to_slv(opcode_type, 16#10#),
      3860 => to_slv(opcode_type, 16#6C#),
      3861 => to_slv(opcode_type, 16#08#),
      3862 => to_slv(opcode_type, 16#06#),
      3863 => to_slv(opcode_type, 16#0C#),
      3864 => to_slv(opcode_type, 16#0D#),
      3865 => to_slv(opcode_type, 16#06#),
      3866 => to_slv(opcode_type, 16#10#),
      3867 => to_slv(opcode_type, 16#36#),
      3868 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#07#),
      3873 => to_slv(opcode_type, 16#07#),
      3874 => to_slv(opcode_type, 16#09#),
      3875 => to_slv(opcode_type, 16#08#),
      3876 => to_slv(opcode_type, 16#0D#),
      3877 => to_slv(opcode_type, 16#11#),
      3878 => to_slv(opcode_type, 16#02#),
      3879 => to_slv(opcode_type, 16#11#),
      3880 => to_slv(opcode_type, 16#06#),
      3881 => to_slv(opcode_type, 16#07#),
      3882 => to_slv(opcode_type, 16#0A#),
      3883 => to_slv(opcode_type, 16#0D#),
      3884 => to_slv(opcode_type, 16#05#),
      3885 => to_slv(opcode_type, 16#0E#),
      3886 => to_slv(opcode_type, 16#09#),
      3887 => to_slv(opcode_type, 16#07#),
      3888 => to_slv(opcode_type, 16#02#),
      3889 => to_slv(opcode_type, 16#0D#),
      3890 => to_slv(opcode_type, 16#08#),
      3891 => to_slv(opcode_type, 16#0E#),
      3892 => to_slv(opcode_type, 16#A3#),
      3893 => to_slv(opcode_type, 16#06#),
      3894 => to_slv(opcode_type, 16#09#),
      3895 => to_slv(opcode_type, 16#60#),
      3896 => to_slv(opcode_type, 16#0A#),
      3897 => to_slv(opcode_type, 16#09#),
      3898 => to_slv(opcode_type, 16#0B#),
      3899 => to_slv(opcode_type, 16#0B#),
      3900 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#06#),
      3905 => to_slv(opcode_type, 16#08#),
      3906 => to_slv(opcode_type, 16#08#),
      3907 => to_slv(opcode_type, 16#08#),
      3908 => to_slv(opcode_type, 16#0F#),
      3909 => to_slv(opcode_type, 16#0F#),
      3910 => to_slv(opcode_type, 16#02#),
      3911 => to_slv(opcode_type, 16#0D#),
      3912 => to_slv(opcode_type, 16#06#),
      3913 => to_slv(opcode_type, 16#07#),
      3914 => to_slv(opcode_type, 16#0A#),
      3915 => to_slv(opcode_type, 16#8C#),
      3916 => to_slv(opcode_type, 16#01#),
      3917 => to_slv(opcode_type, 16#DA#),
      3918 => to_slv(opcode_type, 16#06#),
      3919 => to_slv(opcode_type, 16#08#),
      3920 => to_slv(opcode_type, 16#07#),
      3921 => to_slv(opcode_type, 16#0B#),
      3922 => to_slv(opcode_type, 16#0D#),
      3923 => to_slv(opcode_type, 16#07#),
      3924 => to_slv(opcode_type, 16#10#),
      3925 => to_slv(opcode_type, 16#0C#),
      3926 => to_slv(opcode_type, 16#08#),
      3927 => to_slv(opcode_type, 16#02#),
      3928 => to_slv(opcode_type, 16#BD#),
      3929 => to_slv(opcode_type, 16#07#),
      3930 => to_slv(opcode_type, 16#F8#),
      3931 => to_slv(opcode_type, 16#F2#),
      3932 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#09#),
      3937 => to_slv(opcode_type, 16#06#),
      3938 => to_slv(opcode_type, 16#02#),
      3939 => to_slv(opcode_type, 16#07#),
      3940 => to_slv(opcode_type, 16#0A#),
      3941 => to_slv(opcode_type, 16#10#),
      3942 => to_slv(opcode_type, 16#07#),
      3943 => to_slv(opcode_type, 16#09#),
      3944 => to_slv(opcode_type, 16#0C#),
      3945 => to_slv(opcode_type, 16#0C#),
      3946 => to_slv(opcode_type, 16#07#),
      3947 => to_slv(opcode_type, 16#10#),
      3948 => to_slv(opcode_type, 16#11#),
      3949 => to_slv(opcode_type, 16#09#),
      3950 => to_slv(opcode_type, 16#09#),
      3951 => to_slv(opcode_type, 16#06#),
      3952 => to_slv(opcode_type, 16#0C#),
      3953 => to_slv(opcode_type, 16#10#),
      3954 => to_slv(opcode_type, 16#07#),
      3955 => to_slv(opcode_type, 16#11#),
      3956 => to_slv(opcode_type, 16#0D#),
      3957 => to_slv(opcode_type, 16#07#),
      3958 => to_slv(opcode_type, 16#08#),
      3959 => to_slv(opcode_type, 16#10#),
      3960 => to_slv(opcode_type, 16#2A#),
      3961 => to_slv(opcode_type, 16#09#),
      3962 => to_slv(opcode_type, 16#11#),
      3963 => to_slv(opcode_type, 16#3A#),
      3964 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#09#),
      3969 => to_slv(opcode_type, 16#07#),
      3970 => to_slv(opcode_type, 16#09#),
      3971 => to_slv(opcode_type, 16#03#),
      3972 => to_slv(opcode_type, 16#0B#),
      3973 => to_slv(opcode_type, 16#08#),
      3974 => to_slv(opcode_type, 16#0B#),
      3975 => to_slv(opcode_type, 16#0B#),
      3976 => to_slv(opcode_type, 16#08#),
      3977 => to_slv(opcode_type, 16#02#),
      3978 => to_slv(opcode_type, 16#0A#),
      3979 => to_slv(opcode_type, 16#07#),
      3980 => to_slv(opcode_type, 16#0F#),
      3981 => to_slv(opcode_type, 16#0F#),
      3982 => to_slv(opcode_type, 16#06#),
      3983 => to_slv(opcode_type, 16#09#),
      3984 => to_slv(opcode_type, 16#04#),
      3985 => to_slv(opcode_type, 16#10#),
      3986 => to_slv(opcode_type, 16#08#),
      3987 => to_slv(opcode_type, 16#0F#),
      3988 => to_slv(opcode_type, 16#10#),
      3989 => to_slv(opcode_type, 16#06#),
      3990 => to_slv(opcode_type, 16#09#),
      3991 => to_slv(opcode_type, 16#10#),
      3992 => to_slv(opcode_type, 16#0B#),
      3993 => to_slv(opcode_type, 16#09#),
      3994 => to_slv(opcode_type, 16#10#),
      3995 => to_slv(opcode_type, 16#0E#),
      3996 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#09#),
      4001 => to_slv(opcode_type, 16#07#),
      4002 => to_slv(opcode_type, 16#03#),
      4003 => to_slv(opcode_type, 16#07#),
      4004 => to_slv(opcode_type, 16#0F#),
      4005 => to_slv(opcode_type, 16#0A#),
      4006 => to_slv(opcode_type, 16#09#),
      4007 => to_slv(opcode_type, 16#08#),
      4008 => to_slv(opcode_type, 16#11#),
      4009 => to_slv(opcode_type, 16#0E#),
      4010 => to_slv(opcode_type, 16#09#),
      4011 => to_slv(opcode_type, 16#10#),
      4012 => to_slv(opcode_type, 16#D5#),
      4013 => to_slv(opcode_type, 16#06#),
      4014 => to_slv(opcode_type, 16#07#),
      4015 => to_slv(opcode_type, 16#09#),
      4016 => to_slv(opcode_type, 16#0B#),
      4017 => to_slv(opcode_type, 16#11#),
      4018 => to_slv(opcode_type, 16#06#),
      4019 => to_slv(opcode_type, 16#0B#),
      4020 => to_slv(opcode_type, 16#0A#),
      4021 => to_slv(opcode_type, 16#08#),
      4022 => to_slv(opcode_type, 16#07#),
      4023 => to_slv(opcode_type, 16#0D#),
      4024 => to_slv(opcode_type, 16#FD#),
      4025 => to_slv(opcode_type, 16#08#),
      4026 => to_slv(opcode_type, 16#11#),
      4027 => to_slv(opcode_type, 16#0A#),
      4028 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#08#),
      4033 => to_slv(opcode_type, 16#08#),
      4034 => to_slv(opcode_type, 16#03#),
      4035 => to_slv(opcode_type, 16#08#),
      4036 => to_slv(opcode_type, 16#0F#),
      4037 => to_slv(opcode_type, 16#4E#),
      4038 => to_slv(opcode_type, 16#09#),
      4039 => to_slv(opcode_type, 16#09#),
      4040 => to_slv(opcode_type, 16#0F#),
      4041 => to_slv(opcode_type, 16#0C#),
      4042 => to_slv(opcode_type, 16#08#),
      4043 => to_slv(opcode_type, 16#0B#),
      4044 => to_slv(opcode_type, 16#10#),
      4045 => to_slv(opcode_type, 16#06#),
      4046 => to_slv(opcode_type, 16#07#),
      4047 => to_slv(opcode_type, 16#06#),
      4048 => to_slv(opcode_type, 16#48#),
      4049 => to_slv(opcode_type, 16#11#),
      4050 => to_slv(opcode_type, 16#08#),
      4051 => to_slv(opcode_type, 16#0B#),
      4052 => to_slv(opcode_type, 16#0E#),
      4053 => to_slv(opcode_type, 16#08#),
      4054 => to_slv(opcode_type, 16#09#),
      4055 => to_slv(opcode_type, 16#11#),
      4056 => to_slv(opcode_type, 16#0E#),
      4057 => to_slv(opcode_type, 16#06#),
      4058 => to_slv(opcode_type, 16#0A#),
      4059 => to_slv(opcode_type, 16#0C#),
      4060 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#06#),
      4065 => to_slv(opcode_type, 16#07#),
      4066 => to_slv(opcode_type, 16#09#),
      4067 => to_slv(opcode_type, 16#02#),
      4068 => to_slv(opcode_type, 16#0B#),
      4069 => to_slv(opcode_type, 16#07#),
      4070 => to_slv(opcode_type, 16#0B#),
      4071 => to_slv(opcode_type, 16#11#),
      4072 => to_slv(opcode_type, 16#08#),
      4073 => to_slv(opcode_type, 16#02#),
      4074 => to_slv(opcode_type, 16#0A#),
      4075 => to_slv(opcode_type, 16#02#),
      4076 => to_slv(opcode_type, 16#0D#),
      4077 => to_slv(opcode_type, 16#06#),
      4078 => to_slv(opcode_type, 16#09#),
      4079 => to_slv(opcode_type, 16#08#),
      4080 => to_slv(opcode_type, 16#0B#),
      4081 => to_slv(opcode_type, 16#10#),
      4082 => to_slv(opcode_type, 16#09#),
      4083 => to_slv(opcode_type, 16#0E#),
      4084 => to_slv(opcode_type, 16#0E#),
      4085 => to_slv(opcode_type, 16#07#),
      4086 => to_slv(opcode_type, 16#06#),
      4087 => to_slv(opcode_type, 16#0C#),
      4088 => to_slv(opcode_type, 16#11#),
      4089 => to_slv(opcode_type, 16#07#),
      4090 => to_slv(opcode_type, 16#0B#),
      4091 => to_slv(opcode_type, 16#11#),
      4092 to 4095 => (others => '0')
  ),

    -- Bin `29`...
    28 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#08#),
      1 => to_slv(opcode_type, 16#07#),
      2 => to_slv(opcode_type, 16#07#),
      3 => to_slv(opcode_type, 16#04#),
      4 => to_slv(opcode_type, 16#0F#),
      5 => to_slv(opcode_type, 16#06#),
      6 => to_slv(opcode_type, 16#0E#),
      7 => to_slv(opcode_type, 16#11#),
      8 => to_slv(opcode_type, 16#06#),
      9 => to_slv(opcode_type, 16#06#),
      10 => to_slv(opcode_type, 16#11#),
      11 => to_slv(opcode_type, 16#3D#),
      12 => to_slv(opcode_type, 16#04#),
      13 => to_slv(opcode_type, 16#0C#),
      14 => to_slv(opcode_type, 16#06#),
      15 => to_slv(opcode_type, 16#06#),
      16 => to_slv(opcode_type, 16#07#),
      17 => to_slv(opcode_type, 16#11#),
      18 => to_slv(opcode_type, 16#0A#),
      19 => to_slv(opcode_type, 16#09#),
      20 => to_slv(opcode_type, 16#0A#),
      21 => to_slv(opcode_type, 16#0F#),
      22 => to_slv(opcode_type, 16#09#),
      23 => to_slv(opcode_type, 16#08#),
      24 => to_slv(opcode_type, 16#0A#),
      25 => to_slv(opcode_type, 16#21#),
      26 => to_slv(opcode_type, 16#06#),
      27 => to_slv(opcode_type, 16#0F#),
      28 => to_slv(opcode_type, 16#0C#),
      29 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#08#),
      33 => to_slv(opcode_type, 16#09#),
      34 => to_slv(opcode_type, 16#08#),
      35 => to_slv(opcode_type, 16#06#),
      36 => to_slv(opcode_type, 16#10#),
      37 => to_slv(opcode_type, 16#0E#),
      38 => to_slv(opcode_type, 16#01#),
      39 => to_slv(opcode_type, 16#0C#),
      40 => to_slv(opcode_type, 16#09#),
      41 => to_slv(opcode_type, 16#02#),
      42 => to_slv(opcode_type, 16#0D#),
      43 => to_slv(opcode_type, 16#08#),
      44 => to_slv(opcode_type, 16#10#),
      45 => to_slv(opcode_type, 16#0E#),
      46 => to_slv(opcode_type, 16#09#),
      47 => to_slv(opcode_type, 16#07#),
      48 => to_slv(opcode_type, 16#09#),
      49 => to_slv(opcode_type, 16#0B#),
      50 => to_slv(opcode_type, 16#0D#),
      51 => to_slv(opcode_type, 16#09#),
      52 => to_slv(opcode_type, 16#0A#),
      53 => to_slv(opcode_type, 16#0E#),
      54 => to_slv(opcode_type, 16#06#),
      55 => to_slv(opcode_type, 16#08#),
      56 => to_slv(opcode_type, 16#2C#),
      57 => to_slv(opcode_type, 16#0F#),
      58 => to_slv(opcode_type, 16#06#),
      59 => to_slv(opcode_type, 16#0C#),
      60 => to_slv(opcode_type, 16#0F#),
      61 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#06#),
      65 => to_slv(opcode_type, 16#09#),
      66 => to_slv(opcode_type, 16#08#),
      67 => to_slv(opcode_type, 16#06#),
      68 => to_slv(opcode_type, 16#0D#),
      69 => to_slv(opcode_type, 16#0D#),
      70 => to_slv(opcode_type, 16#07#),
      71 => to_slv(opcode_type, 16#0D#),
      72 => to_slv(opcode_type, 16#32#),
      73 => to_slv(opcode_type, 16#07#),
      74 => to_slv(opcode_type, 16#03#),
      75 => to_slv(opcode_type, 16#0C#),
      76 => to_slv(opcode_type, 16#01#),
      77 => to_slv(opcode_type, 16#0E#),
      78 => to_slv(opcode_type, 16#07#),
      79 => to_slv(opcode_type, 16#07#),
      80 => to_slv(opcode_type, 16#06#),
      81 => to_slv(opcode_type, 16#11#),
      82 => to_slv(opcode_type, 16#0D#),
      83 => to_slv(opcode_type, 16#07#),
      84 => to_slv(opcode_type, 16#0D#),
      85 => to_slv(opcode_type, 16#0A#),
      86 => to_slv(opcode_type, 16#07#),
      87 => to_slv(opcode_type, 16#08#),
      88 => to_slv(opcode_type, 16#0C#),
      89 => to_slv(opcode_type, 16#0B#),
      90 => to_slv(opcode_type, 16#06#),
      91 => to_slv(opcode_type, 16#0C#),
      92 => to_slv(opcode_type, 16#55#),
      93 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#08#),
      97 => to_slv(opcode_type, 16#09#),
      98 => to_slv(opcode_type, 16#07#),
      99 => to_slv(opcode_type, 16#08#),
      100 => to_slv(opcode_type, 16#0F#),
      101 => to_slv(opcode_type, 16#11#),
      102 => to_slv(opcode_type, 16#01#),
      103 => to_slv(opcode_type, 16#11#),
      104 => to_slv(opcode_type, 16#07#),
      105 => to_slv(opcode_type, 16#04#),
      106 => to_slv(opcode_type, 16#0B#),
      107 => to_slv(opcode_type, 16#06#),
      108 => to_slv(opcode_type, 16#0A#),
      109 => to_slv(opcode_type, 16#11#),
      110 => to_slv(opcode_type, 16#07#),
      111 => to_slv(opcode_type, 16#08#),
      112 => to_slv(opcode_type, 16#07#),
      113 => to_slv(opcode_type, 16#0C#),
      114 => to_slv(opcode_type, 16#11#),
      115 => to_slv(opcode_type, 16#08#),
      116 => to_slv(opcode_type, 16#11#),
      117 => to_slv(opcode_type, 16#0E#),
      118 => to_slv(opcode_type, 16#06#),
      119 => to_slv(opcode_type, 16#09#),
      120 => to_slv(opcode_type, 16#0F#),
      121 => to_slv(opcode_type, 16#0B#),
      122 => to_slv(opcode_type, 16#08#),
      123 => to_slv(opcode_type, 16#0D#),
      124 => to_slv(opcode_type, 16#0D#),
      125 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#07#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#06#),
      131 => to_slv(opcode_type, 16#02#),
      132 => to_slv(opcode_type, 16#0E#),
      133 => to_slv(opcode_type, 16#03#),
      134 => to_slv(opcode_type, 16#0A#),
      135 => to_slv(opcode_type, 16#06#),
      136 => to_slv(opcode_type, 16#06#),
      137 => to_slv(opcode_type, 16#11#),
      138 => to_slv(opcode_type, 16#10#),
      139 => to_slv(opcode_type, 16#09#),
      140 => to_slv(opcode_type, 16#10#),
      141 => to_slv(opcode_type, 16#0F#),
      142 => to_slv(opcode_type, 16#07#),
      143 => to_slv(opcode_type, 16#09#),
      144 => to_slv(opcode_type, 16#09#),
      145 => to_slv(opcode_type, 16#0E#),
      146 => to_slv(opcode_type, 16#0D#),
      147 => to_slv(opcode_type, 16#07#),
      148 => to_slv(opcode_type, 16#0E#),
      149 => to_slv(opcode_type, 16#0C#),
      150 => to_slv(opcode_type, 16#06#),
      151 => to_slv(opcode_type, 16#08#),
      152 => to_slv(opcode_type, 16#1F#),
      153 => to_slv(opcode_type, 16#10#),
      154 => to_slv(opcode_type, 16#08#),
      155 => to_slv(opcode_type, 16#0C#),
      156 => to_slv(opcode_type, 16#0F#),
      157 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#08#),
      161 => to_slv(opcode_type, 16#07#),
      162 => to_slv(opcode_type, 16#08#),
      163 => to_slv(opcode_type, 16#05#),
      164 => to_slv(opcode_type, 16#0C#),
      165 => to_slv(opcode_type, 16#02#),
      166 => to_slv(opcode_type, 16#10#),
      167 => to_slv(opcode_type, 16#08#),
      168 => to_slv(opcode_type, 16#09#),
      169 => to_slv(opcode_type, 16#0E#),
      170 => to_slv(opcode_type, 16#0C#),
      171 => to_slv(opcode_type, 16#07#),
      172 => to_slv(opcode_type, 16#0D#),
      173 => to_slv(opcode_type, 16#0C#),
      174 => to_slv(opcode_type, 16#09#),
      175 => to_slv(opcode_type, 16#07#),
      176 => to_slv(opcode_type, 16#08#),
      177 => to_slv(opcode_type, 16#0B#),
      178 => to_slv(opcode_type, 16#0D#),
      179 => to_slv(opcode_type, 16#07#),
      180 => to_slv(opcode_type, 16#6D#),
      181 => to_slv(opcode_type, 16#0D#),
      182 => to_slv(opcode_type, 16#09#),
      183 => to_slv(opcode_type, 16#09#),
      184 => to_slv(opcode_type, 16#0C#),
      185 => to_slv(opcode_type, 16#0A#),
      186 => to_slv(opcode_type, 16#07#),
      187 => to_slv(opcode_type, 16#0B#),
      188 => to_slv(opcode_type, 16#0E#),
      189 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#08#),
      193 => to_slv(opcode_type, 16#06#),
      194 => to_slv(opcode_type, 16#09#),
      195 => to_slv(opcode_type, 16#02#),
      196 => to_slv(opcode_type, 16#10#),
      197 => to_slv(opcode_type, 16#03#),
      198 => to_slv(opcode_type, 16#49#),
      199 => to_slv(opcode_type, 16#09#),
      200 => to_slv(opcode_type, 16#09#),
      201 => to_slv(opcode_type, 16#0E#),
      202 => to_slv(opcode_type, 16#10#),
      203 => to_slv(opcode_type, 16#09#),
      204 => to_slv(opcode_type, 16#0F#),
      205 => to_slv(opcode_type, 16#0B#),
      206 => to_slv(opcode_type, 16#07#),
      207 => to_slv(opcode_type, 16#08#),
      208 => to_slv(opcode_type, 16#06#),
      209 => to_slv(opcode_type, 16#0E#),
      210 => to_slv(opcode_type, 16#0C#),
      211 => to_slv(opcode_type, 16#06#),
      212 => to_slv(opcode_type, 16#0D#),
      213 => to_slv(opcode_type, 16#0F#),
      214 => to_slv(opcode_type, 16#07#),
      215 => to_slv(opcode_type, 16#09#),
      216 => to_slv(opcode_type, 16#0A#),
      217 => to_slv(opcode_type, 16#0B#),
      218 => to_slv(opcode_type, 16#09#),
      219 => to_slv(opcode_type, 16#10#),
      220 => to_slv(opcode_type, 16#0E#),
      221 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#09#),
      225 => to_slv(opcode_type, 16#09#),
      226 => to_slv(opcode_type, 16#06#),
      227 => to_slv(opcode_type, 16#03#),
      228 => to_slv(opcode_type, 16#0D#),
      229 => to_slv(opcode_type, 16#03#),
      230 => to_slv(opcode_type, 16#0E#),
      231 => to_slv(opcode_type, 16#07#),
      232 => to_slv(opcode_type, 16#09#),
      233 => to_slv(opcode_type, 16#0C#),
      234 => to_slv(opcode_type, 16#0D#),
      235 => to_slv(opcode_type, 16#06#),
      236 => to_slv(opcode_type, 16#11#),
      237 => to_slv(opcode_type, 16#0E#),
      238 => to_slv(opcode_type, 16#06#),
      239 => to_slv(opcode_type, 16#09#),
      240 => to_slv(opcode_type, 16#07#),
      241 => to_slv(opcode_type, 16#10#),
      242 => to_slv(opcode_type, 16#0B#),
      243 => to_slv(opcode_type, 16#09#),
      244 => to_slv(opcode_type, 16#0B#),
      245 => to_slv(opcode_type, 16#47#),
      246 => to_slv(opcode_type, 16#08#),
      247 => to_slv(opcode_type, 16#08#),
      248 => to_slv(opcode_type, 16#0A#),
      249 => to_slv(opcode_type, 16#0B#),
      250 => to_slv(opcode_type, 16#09#),
      251 => to_slv(opcode_type, 16#0D#),
      252 => to_slv(opcode_type, 16#10#),
      253 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#07#),
      257 => to_slv(opcode_type, 16#09#),
      258 => to_slv(opcode_type, 16#09#),
      259 => to_slv(opcode_type, 16#06#),
      260 => to_slv(opcode_type, 16#A1#),
      261 => to_slv(opcode_type, 16#0E#),
      262 => to_slv(opcode_type, 16#05#),
      263 => to_slv(opcode_type, 16#0C#),
      264 => to_slv(opcode_type, 16#07#),
      265 => to_slv(opcode_type, 16#06#),
      266 => to_slv(opcode_type, 16#0C#),
      267 => to_slv(opcode_type, 16#0C#),
      268 => to_slv(opcode_type, 16#03#),
      269 => to_slv(opcode_type, 16#0C#),
      270 => to_slv(opcode_type, 16#06#),
      271 => to_slv(opcode_type, 16#06#),
      272 => to_slv(opcode_type, 16#08#),
      273 => to_slv(opcode_type, 16#10#),
      274 => to_slv(opcode_type, 16#11#),
      275 => to_slv(opcode_type, 16#07#),
      276 => to_slv(opcode_type, 16#11#),
      277 => to_slv(opcode_type, 16#0F#),
      278 => to_slv(opcode_type, 16#07#),
      279 => to_slv(opcode_type, 16#08#),
      280 => to_slv(opcode_type, 16#0A#),
      281 => to_slv(opcode_type, 16#10#),
      282 => to_slv(opcode_type, 16#06#),
      283 => to_slv(opcode_type, 16#0E#),
      284 => to_slv(opcode_type, 16#0E#),
      285 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#06#),
      289 => to_slv(opcode_type, 16#07#),
      290 => to_slv(opcode_type, 16#07#),
      291 => to_slv(opcode_type, 16#06#),
      292 => to_slv(opcode_type, 16#0A#),
      293 => to_slv(opcode_type, 16#0F#),
      294 => to_slv(opcode_type, 16#01#),
      295 => to_slv(opcode_type, 16#0A#),
      296 => to_slv(opcode_type, 16#08#),
      297 => to_slv(opcode_type, 16#04#),
      298 => to_slv(opcode_type, 16#11#),
      299 => to_slv(opcode_type, 16#06#),
      300 => to_slv(opcode_type, 16#0B#),
      301 => to_slv(opcode_type, 16#10#),
      302 => to_slv(opcode_type, 16#08#),
      303 => to_slv(opcode_type, 16#06#),
      304 => to_slv(opcode_type, 16#09#),
      305 => to_slv(opcode_type, 16#0D#),
      306 => to_slv(opcode_type, 16#10#),
      307 => to_slv(opcode_type, 16#06#),
      308 => to_slv(opcode_type, 16#0A#),
      309 => to_slv(opcode_type, 16#0C#),
      310 => to_slv(opcode_type, 16#08#),
      311 => to_slv(opcode_type, 16#07#),
      312 => to_slv(opcode_type, 16#11#),
      313 => to_slv(opcode_type, 16#0A#),
      314 => to_slv(opcode_type, 16#07#),
      315 => to_slv(opcode_type, 16#0F#),
      316 => to_slv(opcode_type, 16#0E#),
      317 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#08#),
      321 => to_slv(opcode_type, 16#08#),
      322 => to_slv(opcode_type, 16#08#),
      323 => to_slv(opcode_type, 16#05#),
      324 => to_slv(opcode_type, 16#0E#),
      325 => to_slv(opcode_type, 16#07#),
      326 => to_slv(opcode_type, 16#0A#),
      327 => to_slv(opcode_type, 16#0F#),
      328 => to_slv(opcode_type, 16#09#),
      329 => to_slv(opcode_type, 16#02#),
      330 => to_slv(opcode_type, 16#0A#),
      331 => to_slv(opcode_type, 16#08#),
      332 => to_slv(opcode_type, 16#0D#),
      333 => to_slv(opcode_type, 16#0F#),
      334 => to_slv(opcode_type, 16#07#),
      335 => to_slv(opcode_type, 16#06#),
      336 => to_slv(opcode_type, 16#07#),
      337 => to_slv(opcode_type, 16#0F#),
      338 => to_slv(opcode_type, 16#0B#),
      339 => to_slv(opcode_type, 16#07#),
      340 => to_slv(opcode_type, 16#0C#),
      341 => to_slv(opcode_type, 16#0F#),
      342 => to_slv(opcode_type, 16#07#),
      343 => to_slv(opcode_type, 16#08#),
      344 => to_slv(opcode_type, 16#B2#),
      345 => to_slv(opcode_type, 16#0E#),
      346 => to_slv(opcode_type, 16#09#),
      347 => to_slv(opcode_type, 16#11#),
      348 => to_slv(opcode_type, 16#0C#),
      349 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#07#),
      353 => to_slv(opcode_type, 16#08#),
      354 => to_slv(opcode_type, 16#07#),
      355 => to_slv(opcode_type, 16#05#),
      356 => to_slv(opcode_type, 16#0F#),
      357 => to_slv(opcode_type, 16#06#),
      358 => to_slv(opcode_type, 16#0B#),
      359 => to_slv(opcode_type, 16#0C#),
      360 => to_slv(opcode_type, 16#06#),
      361 => to_slv(opcode_type, 16#08#),
      362 => to_slv(opcode_type, 16#0E#),
      363 => to_slv(opcode_type, 16#0F#),
      364 => to_slv(opcode_type, 16#04#),
      365 => to_slv(opcode_type, 16#0D#),
      366 => to_slv(opcode_type, 16#07#),
      367 => to_slv(opcode_type, 16#09#),
      368 => to_slv(opcode_type, 16#09#),
      369 => to_slv(opcode_type, 16#0D#),
      370 => to_slv(opcode_type, 16#0E#),
      371 => to_slv(opcode_type, 16#09#),
      372 => to_slv(opcode_type, 16#96#),
      373 => to_slv(opcode_type, 16#0A#),
      374 => to_slv(opcode_type, 16#07#),
      375 => to_slv(opcode_type, 16#09#),
      376 => to_slv(opcode_type, 16#A1#),
      377 => to_slv(opcode_type, 16#0F#),
      378 => to_slv(opcode_type, 16#06#),
      379 => to_slv(opcode_type, 16#0B#),
      380 => to_slv(opcode_type, 16#11#),
      381 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#09#),
      385 => to_slv(opcode_type, 16#06#),
      386 => to_slv(opcode_type, 16#07#),
      387 => to_slv(opcode_type, 16#03#),
      388 => to_slv(opcode_type, 16#0D#),
      389 => to_slv(opcode_type, 16#07#),
      390 => to_slv(opcode_type, 16#10#),
      391 => to_slv(opcode_type, 16#0C#),
      392 => to_slv(opcode_type, 16#06#),
      393 => to_slv(opcode_type, 16#04#),
      394 => to_slv(opcode_type, 16#0D#),
      395 => to_slv(opcode_type, 16#07#),
      396 => to_slv(opcode_type, 16#0B#),
      397 => to_slv(opcode_type, 16#0D#),
      398 => to_slv(opcode_type, 16#08#),
      399 => to_slv(opcode_type, 16#08#),
      400 => to_slv(opcode_type, 16#06#),
      401 => to_slv(opcode_type, 16#0E#),
      402 => to_slv(opcode_type, 16#0E#),
      403 => to_slv(opcode_type, 16#08#),
      404 => to_slv(opcode_type, 16#11#),
      405 => to_slv(opcode_type, 16#0F#),
      406 => to_slv(opcode_type, 16#09#),
      407 => to_slv(opcode_type, 16#07#),
      408 => to_slv(opcode_type, 16#11#),
      409 => to_slv(opcode_type, 16#0F#),
      410 => to_slv(opcode_type, 16#09#),
      411 => to_slv(opcode_type, 16#0A#),
      412 => to_slv(opcode_type, 16#0E#),
      413 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#09#),
      417 => to_slv(opcode_type, 16#06#),
      418 => to_slv(opcode_type, 16#06#),
      419 => to_slv(opcode_type, 16#05#),
      420 => to_slv(opcode_type, 16#0A#),
      421 => to_slv(opcode_type, 16#02#),
      422 => to_slv(opcode_type, 16#10#),
      423 => to_slv(opcode_type, 16#06#),
      424 => to_slv(opcode_type, 16#07#),
      425 => to_slv(opcode_type, 16#0C#),
      426 => to_slv(opcode_type, 16#0F#),
      427 => to_slv(opcode_type, 16#08#),
      428 => to_slv(opcode_type, 16#0F#),
      429 => to_slv(opcode_type, 16#0C#),
      430 => to_slv(opcode_type, 16#06#),
      431 => to_slv(opcode_type, 16#06#),
      432 => to_slv(opcode_type, 16#06#),
      433 => to_slv(opcode_type, 16#0E#),
      434 => to_slv(opcode_type, 16#11#),
      435 => to_slv(opcode_type, 16#07#),
      436 => to_slv(opcode_type, 16#10#),
      437 => to_slv(opcode_type, 16#0E#),
      438 => to_slv(opcode_type, 16#06#),
      439 => to_slv(opcode_type, 16#07#),
      440 => to_slv(opcode_type, 16#0D#),
      441 => to_slv(opcode_type, 16#0B#),
      442 => to_slv(opcode_type, 16#09#),
      443 => to_slv(opcode_type, 16#0D#),
      444 => to_slv(opcode_type, 16#11#),
      445 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#07#),
      449 => to_slv(opcode_type, 16#06#),
      450 => to_slv(opcode_type, 16#08#),
      451 => to_slv(opcode_type, 16#06#),
      452 => to_slv(opcode_type, 16#0A#),
      453 => to_slv(opcode_type, 16#0D#),
      454 => to_slv(opcode_type, 16#05#),
      455 => to_slv(opcode_type, 16#0B#),
      456 => to_slv(opcode_type, 16#08#),
      457 => to_slv(opcode_type, 16#04#),
      458 => to_slv(opcode_type, 16#0F#),
      459 => to_slv(opcode_type, 16#06#),
      460 => to_slv(opcode_type, 16#11#),
      461 => to_slv(opcode_type, 16#0B#),
      462 => to_slv(opcode_type, 16#09#),
      463 => to_slv(opcode_type, 16#09#),
      464 => to_slv(opcode_type, 16#07#),
      465 => to_slv(opcode_type, 16#99#),
      466 => to_slv(opcode_type, 16#0A#),
      467 => to_slv(opcode_type, 16#08#),
      468 => to_slv(opcode_type, 16#0E#),
      469 => to_slv(opcode_type, 16#7B#),
      470 => to_slv(opcode_type, 16#07#),
      471 => to_slv(opcode_type, 16#07#),
      472 => to_slv(opcode_type, 16#0B#),
      473 => to_slv(opcode_type, 16#0D#),
      474 => to_slv(opcode_type, 16#06#),
      475 => to_slv(opcode_type, 16#0F#),
      476 => to_slv(opcode_type, 16#0B#),
      477 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#07#),
      481 => to_slv(opcode_type, 16#07#),
      482 => to_slv(opcode_type, 16#09#),
      483 => to_slv(opcode_type, 16#07#),
      484 => to_slv(opcode_type, 16#0F#),
      485 => to_slv(opcode_type, 16#10#),
      486 => to_slv(opcode_type, 16#05#),
      487 => to_slv(opcode_type, 16#0E#),
      488 => to_slv(opcode_type, 16#06#),
      489 => to_slv(opcode_type, 16#03#),
      490 => to_slv(opcode_type, 16#10#),
      491 => to_slv(opcode_type, 16#08#),
      492 => to_slv(opcode_type, 16#0D#),
      493 => to_slv(opcode_type, 16#10#),
      494 => to_slv(opcode_type, 16#08#),
      495 => to_slv(opcode_type, 16#08#),
      496 => to_slv(opcode_type, 16#09#),
      497 => to_slv(opcode_type, 16#0E#),
      498 => to_slv(opcode_type, 16#ED#),
      499 => to_slv(opcode_type, 16#09#),
      500 => to_slv(opcode_type, 16#0A#),
      501 => to_slv(opcode_type, 16#0C#),
      502 => to_slv(opcode_type, 16#06#),
      503 => to_slv(opcode_type, 16#07#),
      504 => to_slv(opcode_type, 16#10#),
      505 => to_slv(opcode_type, 16#0E#),
      506 => to_slv(opcode_type, 16#08#),
      507 => to_slv(opcode_type, 16#0F#),
      508 => to_slv(opcode_type, 16#0C#),
      509 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#06#),
      514 => to_slv(opcode_type, 16#08#),
      515 => to_slv(opcode_type, 16#05#),
      516 => to_slv(opcode_type, 16#10#),
      517 => to_slv(opcode_type, 16#07#),
      518 => to_slv(opcode_type, 16#0D#),
      519 => to_slv(opcode_type, 16#1C#),
      520 => to_slv(opcode_type, 16#08#),
      521 => to_slv(opcode_type, 16#01#),
      522 => to_slv(opcode_type, 16#0C#),
      523 => to_slv(opcode_type, 16#08#),
      524 => to_slv(opcode_type, 16#0C#),
      525 => to_slv(opcode_type, 16#0A#),
      526 => to_slv(opcode_type, 16#07#),
      527 => to_slv(opcode_type, 16#06#),
      528 => to_slv(opcode_type, 16#07#),
      529 => to_slv(opcode_type, 16#11#),
      530 => to_slv(opcode_type, 16#0F#),
      531 => to_slv(opcode_type, 16#09#),
      532 => to_slv(opcode_type, 16#0D#),
      533 => to_slv(opcode_type, 16#1D#),
      534 => to_slv(opcode_type, 16#08#),
      535 => to_slv(opcode_type, 16#09#),
      536 => to_slv(opcode_type, 16#10#),
      537 => to_slv(opcode_type, 16#0A#),
      538 => to_slv(opcode_type, 16#08#),
      539 => to_slv(opcode_type, 16#0B#),
      540 => to_slv(opcode_type, 16#0D#),
      541 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#07#),
      545 => to_slv(opcode_type, 16#08#),
      546 => to_slv(opcode_type, 16#06#),
      547 => to_slv(opcode_type, 16#01#),
      548 => to_slv(opcode_type, 16#0F#),
      549 => to_slv(opcode_type, 16#02#),
      550 => to_slv(opcode_type, 16#0F#),
      551 => to_slv(opcode_type, 16#06#),
      552 => to_slv(opcode_type, 16#08#),
      553 => to_slv(opcode_type, 16#0B#),
      554 => to_slv(opcode_type, 16#0A#),
      555 => to_slv(opcode_type, 16#08#),
      556 => to_slv(opcode_type, 16#0D#),
      557 => to_slv(opcode_type, 16#0B#),
      558 => to_slv(opcode_type, 16#09#),
      559 => to_slv(opcode_type, 16#06#),
      560 => to_slv(opcode_type, 16#08#),
      561 => to_slv(opcode_type, 16#10#),
      562 => to_slv(opcode_type, 16#0E#),
      563 => to_slv(opcode_type, 16#06#),
      564 => to_slv(opcode_type, 16#11#),
      565 => to_slv(opcode_type, 16#0E#),
      566 => to_slv(opcode_type, 16#09#),
      567 => to_slv(opcode_type, 16#09#),
      568 => to_slv(opcode_type, 16#0B#),
      569 => to_slv(opcode_type, 16#0E#),
      570 => to_slv(opcode_type, 16#09#),
      571 => to_slv(opcode_type, 16#10#),
      572 => to_slv(opcode_type, 16#10#),
      573 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#08#),
      577 => to_slv(opcode_type, 16#09#),
      578 => to_slv(opcode_type, 16#09#),
      579 => to_slv(opcode_type, 16#04#),
      580 => to_slv(opcode_type, 16#0D#),
      581 => to_slv(opcode_type, 16#05#),
      582 => to_slv(opcode_type, 16#10#),
      583 => to_slv(opcode_type, 16#09#),
      584 => to_slv(opcode_type, 16#09#),
      585 => to_slv(opcode_type, 16#11#),
      586 => to_slv(opcode_type, 16#0A#),
      587 => to_slv(opcode_type, 16#08#),
      588 => to_slv(opcode_type, 16#0D#),
      589 => to_slv(opcode_type, 16#0F#),
      590 => to_slv(opcode_type, 16#08#),
      591 => to_slv(opcode_type, 16#07#),
      592 => to_slv(opcode_type, 16#08#),
      593 => to_slv(opcode_type, 16#11#),
      594 => to_slv(opcode_type, 16#0C#),
      595 => to_slv(opcode_type, 16#07#),
      596 => to_slv(opcode_type, 16#7E#),
      597 => to_slv(opcode_type, 16#0D#),
      598 => to_slv(opcode_type, 16#07#),
      599 => to_slv(opcode_type, 16#07#),
      600 => to_slv(opcode_type, 16#11#),
      601 => to_slv(opcode_type, 16#0F#),
      602 => to_slv(opcode_type, 16#08#),
      603 => to_slv(opcode_type, 16#0B#),
      604 => to_slv(opcode_type, 16#0C#),
      605 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#08#),
      609 => to_slv(opcode_type, 16#07#),
      610 => to_slv(opcode_type, 16#09#),
      611 => to_slv(opcode_type, 16#03#),
      612 => to_slv(opcode_type, 16#0A#),
      613 => to_slv(opcode_type, 16#07#),
      614 => to_slv(opcode_type, 16#11#),
      615 => to_slv(opcode_type, 16#0A#),
      616 => to_slv(opcode_type, 16#08#),
      617 => to_slv(opcode_type, 16#02#),
      618 => to_slv(opcode_type, 16#78#),
      619 => to_slv(opcode_type, 16#07#),
      620 => to_slv(opcode_type, 16#0E#),
      621 => to_slv(opcode_type, 16#10#),
      622 => to_slv(opcode_type, 16#06#),
      623 => to_slv(opcode_type, 16#06#),
      624 => to_slv(opcode_type, 16#07#),
      625 => to_slv(opcode_type, 16#0D#),
      626 => to_slv(opcode_type, 16#11#),
      627 => to_slv(opcode_type, 16#09#),
      628 => to_slv(opcode_type, 16#11#),
      629 => to_slv(opcode_type, 16#0F#),
      630 => to_slv(opcode_type, 16#08#),
      631 => to_slv(opcode_type, 16#08#),
      632 => to_slv(opcode_type, 16#10#),
      633 => to_slv(opcode_type, 16#DD#),
      634 => to_slv(opcode_type, 16#08#),
      635 => to_slv(opcode_type, 16#0B#),
      636 => to_slv(opcode_type, 16#88#),
      637 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#06#),
      641 => to_slv(opcode_type, 16#08#),
      642 => to_slv(opcode_type, 16#07#),
      643 => to_slv(opcode_type, 16#02#),
      644 => to_slv(opcode_type, 16#0E#),
      645 => to_slv(opcode_type, 16#04#),
      646 => to_slv(opcode_type, 16#0B#),
      647 => to_slv(opcode_type, 16#06#),
      648 => to_slv(opcode_type, 16#08#),
      649 => to_slv(opcode_type, 16#0B#),
      650 => to_slv(opcode_type, 16#3F#),
      651 => to_slv(opcode_type, 16#07#),
      652 => to_slv(opcode_type, 16#0D#),
      653 => to_slv(opcode_type, 16#0B#),
      654 => to_slv(opcode_type, 16#09#),
      655 => to_slv(opcode_type, 16#06#),
      656 => to_slv(opcode_type, 16#07#),
      657 => to_slv(opcode_type, 16#0B#),
      658 => to_slv(opcode_type, 16#0A#),
      659 => to_slv(opcode_type, 16#08#),
      660 => to_slv(opcode_type, 16#43#),
      661 => to_slv(opcode_type, 16#11#),
      662 => to_slv(opcode_type, 16#07#),
      663 => to_slv(opcode_type, 16#09#),
      664 => to_slv(opcode_type, 16#0B#),
      665 => to_slv(opcode_type, 16#0B#),
      666 => to_slv(opcode_type, 16#08#),
      667 => to_slv(opcode_type, 16#0A#),
      668 => to_slv(opcode_type, 16#0B#),
      669 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#07#),
      673 => to_slv(opcode_type, 16#07#),
      674 => to_slv(opcode_type, 16#07#),
      675 => to_slv(opcode_type, 16#09#),
      676 => to_slv(opcode_type, 16#0E#),
      677 => to_slv(opcode_type, 16#0F#),
      678 => to_slv(opcode_type, 16#09#),
      679 => to_slv(opcode_type, 16#0C#),
      680 => to_slv(opcode_type, 16#0E#),
      681 => to_slv(opcode_type, 16#06#),
      682 => to_slv(opcode_type, 16#05#),
      683 => to_slv(opcode_type, 16#0F#),
      684 => to_slv(opcode_type, 16#02#),
      685 => to_slv(opcode_type, 16#EA#),
      686 => to_slv(opcode_type, 16#07#),
      687 => to_slv(opcode_type, 16#07#),
      688 => to_slv(opcode_type, 16#06#),
      689 => to_slv(opcode_type, 16#0B#),
      690 => to_slv(opcode_type, 16#0C#),
      691 => to_slv(opcode_type, 16#06#),
      692 => to_slv(opcode_type, 16#21#),
      693 => to_slv(opcode_type, 16#11#),
      694 => to_slv(opcode_type, 16#08#),
      695 => to_slv(opcode_type, 16#09#),
      696 => to_slv(opcode_type, 16#24#),
      697 => to_slv(opcode_type, 16#11#),
      698 => to_slv(opcode_type, 16#09#),
      699 => to_slv(opcode_type, 16#64#),
      700 => to_slv(opcode_type, 16#0C#),
      701 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#06#),
      705 => to_slv(opcode_type, 16#08#),
      706 => to_slv(opcode_type, 16#06#),
      707 => to_slv(opcode_type, 16#09#),
      708 => to_slv(opcode_type, 16#0B#),
      709 => to_slv(opcode_type, 16#0F#),
      710 => to_slv(opcode_type, 16#02#),
      711 => to_slv(opcode_type, 16#CB#),
      712 => to_slv(opcode_type, 16#08#),
      713 => to_slv(opcode_type, 16#03#),
      714 => to_slv(opcode_type, 16#11#),
      715 => to_slv(opcode_type, 16#08#),
      716 => to_slv(opcode_type, 16#0F#),
      717 => to_slv(opcode_type, 16#0C#),
      718 => to_slv(opcode_type, 16#07#),
      719 => to_slv(opcode_type, 16#06#),
      720 => to_slv(opcode_type, 16#08#),
      721 => to_slv(opcode_type, 16#10#),
      722 => to_slv(opcode_type, 16#0D#),
      723 => to_slv(opcode_type, 16#06#),
      724 => to_slv(opcode_type, 16#10#),
      725 => to_slv(opcode_type, 16#0A#),
      726 => to_slv(opcode_type, 16#09#),
      727 => to_slv(opcode_type, 16#08#),
      728 => to_slv(opcode_type, 16#10#),
      729 => to_slv(opcode_type, 16#11#),
      730 => to_slv(opcode_type, 16#07#),
      731 => to_slv(opcode_type, 16#0B#),
      732 => to_slv(opcode_type, 16#0E#),
      733 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#07#),
      737 => to_slv(opcode_type, 16#09#),
      738 => to_slv(opcode_type, 16#06#),
      739 => to_slv(opcode_type, 16#09#),
      740 => to_slv(opcode_type, 16#0E#),
      741 => to_slv(opcode_type, 16#0B#),
      742 => to_slv(opcode_type, 16#05#),
      743 => to_slv(opcode_type, 16#E6#),
      744 => to_slv(opcode_type, 16#06#),
      745 => to_slv(opcode_type, 16#05#),
      746 => to_slv(opcode_type, 16#11#),
      747 => to_slv(opcode_type, 16#06#),
      748 => to_slv(opcode_type, 16#0F#),
      749 => to_slv(opcode_type, 16#0D#),
      750 => to_slv(opcode_type, 16#06#),
      751 => to_slv(opcode_type, 16#07#),
      752 => to_slv(opcode_type, 16#08#),
      753 => to_slv(opcode_type, 16#0D#),
      754 => to_slv(opcode_type, 16#0A#),
      755 => to_slv(opcode_type, 16#09#),
      756 => to_slv(opcode_type, 16#0A#),
      757 => to_slv(opcode_type, 16#0C#),
      758 => to_slv(opcode_type, 16#09#),
      759 => to_slv(opcode_type, 16#09#),
      760 => to_slv(opcode_type, 16#0C#),
      761 => to_slv(opcode_type, 16#10#),
      762 => to_slv(opcode_type, 16#09#),
      763 => to_slv(opcode_type, 16#0F#),
      764 => to_slv(opcode_type, 16#10#),
      765 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#06#),
      769 => to_slv(opcode_type, 16#09#),
      770 => to_slv(opcode_type, 16#07#),
      771 => to_slv(opcode_type, 16#05#),
      772 => to_slv(opcode_type, 16#0F#),
      773 => to_slv(opcode_type, 16#03#),
      774 => to_slv(opcode_type, 16#0C#),
      775 => to_slv(opcode_type, 16#08#),
      776 => to_slv(opcode_type, 16#08#),
      777 => to_slv(opcode_type, 16#BE#),
      778 => to_slv(opcode_type, 16#0E#),
      779 => to_slv(opcode_type, 16#06#),
      780 => to_slv(opcode_type, 16#0A#),
      781 => to_slv(opcode_type, 16#0D#),
      782 => to_slv(opcode_type, 16#09#),
      783 => to_slv(opcode_type, 16#09#),
      784 => to_slv(opcode_type, 16#08#),
      785 => to_slv(opcode_type, 16#10#),
      786 => to_slv(opcode_type, 16#12#),
      787 => to_slv(opcode_type, 16#08#),
      788 => to_slv(opcode_type, 16#36#),
      789 => to_slv(opcode_type, 16#0E#),
      790 => to_slv(opcode_type, 16#07#),
      791 => to_slv(opcode_type, 16#07#),
      792 => to_slv(opcode_type, 16#10#),
      793 => to_slv(opcode_type, 16#10#),
      794 => to_slv(opcode_type, 16#09#),
      795 => to_slv(opcode_type, 16#0B#),
      796 => to_slv(opcode_type, 16#0A#),
      797 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#08#),
      801 => to_slv(opcode_type, 16#08#),
      802 => to_slv(opcode_type, 16#07#),
      803 => to_slv(opcode_type, 16#03#),
      804 => to_slv(opcode_type, 16#0B#),
      805 => to_slv(opcode_type, 16#02#),
      806 => to_slv(opcode_type, 16#0B#),
      807 => to_slv(opcode_type, 16#08#),
      808 => to_slv(opcode_type, 16#07#),
      809 => to_slv(opcode_type, 16#0B#),
      810 => to_slv(opcode_type, 16#10#),
      811 => to_slv(opcode_type, 16#08#),
      812 => to_slv(opcode_type, 16#0A#),
      813 => to_slv(opcode_type, 16#0B#),
      814 => to_slv(opcode_type, 16#06#),
      815 => to_slv(opcode_type, 16#06#),
      816 => to_slv(opcode_type, 16#09#),
      817 => to_slv(opcode_type, 16#10#),
      818 => to_slv(opcode_type, 16#0F#),
      819 => to_slv(opcode_type, 16#09#),
      820 => to_slv(opcode_type, 16#0D#),
      821 => to_slv(opcode_type, 16#0B#),
      822 => to_slv(opcode_type, 16#07#),
      823 => to_slv(opcode_type, 16#09#),
      824 => to_slv(opcode_type, 16#0C#),
      825 => to_slv(opcode_type, 16#0A#),
      826 => to_slv(opcode_type, 16#06#),
      827 => to_slv(opcode_type, 16#FF#),
      828 => to_slv(opcode_type, 16#0E#),
      829 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#08#),
      833 => to_slv(opcode_type, 16#06#),
      834 => to_slv(opcode_type, 16#09#),
      835 => to_slv(opcode_type, 16#06#),
      836 => to_slv(opcode_type, 16#78#),
      837 => to_slv(opcode_type, 16#0A#),
      838 => to_slv(opcode_type, 16#08#),
      839 => to_slv(opcode_type, 16#CD#),
      840 => to_slv(opcode_type, 16#0B#),
      841 => to_slv(opcode_type, 16#08#),
      842 => to_slv(opcode_type, 16#05#),
      843 => to_slv(opcode_type, 16#B8#),
      844 => to_slv(opcode_type, 16#03#),
      845 => to_slv(opcode_type, 16#11#),
      846 => to_slv(opcode_type, 16#08#),
      847 => to_slv(opcode_type, 16#08#),
      848 => to_slv(opcode_type, 16#07#),
      849 => to_slv(opcode_type, 16#0D#),
      850 => to_slv(opcode_type, 16#0A#),
      851 => to_slv(opcode_type, 16#07#),
      852 => to_slv(opcode_type, 16#10#),
      853 => to_slv(opcode_type, 16#0F#),
      854 => to_slv(opcode_type, 16#06#),
      855 => to_slv(opcode_type, 16#07#),
      856 => to_slv(opcode_type, 16#10#),
      857 => to_slv(opcode_type, 16#10#),
      858 => to_slv(opcode_type, 16#09#),
      859 => to_slv(opcode_type, 16#0A#),
      860 => to_slv(opcode_type, 16#0F#),
      861 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#07#),
      865 => to_slv(opcode_type, 16#07#),
      866 => to_slv(opcode_type, 16#09#),
      867 => to_slv(opcode_type, 16#08#),
      868 => to_slv(opcode_type, 16#10#),
      869 => to_slv(opcode_type, 16#0F#),
      870 => to_slv(opcode_type, 16#07#),
      871 => to_slv(opcode_type, 16#0B#),
      872 => to_slv(opcode_type, 16#EC#),
      873 => to_slv(opcode_type, 16#09#),
      874 => to_slv(opcode_type, 16#06#),
      875 => to_slv(opcode_type, 16#0E#),
      876 => to_slv(opcode_type, 16#11#),
      877 => to_slv(opcode_type, 16#06#),
      878 => to_slv(opcode_type, 16#0F#),
      879 => to_slv(opcode_type, 16#10#),
      880 => to_slv(opcode_type, 16#06#),
      881 => to_slv(opcode_type, 16#07#),
      882 => to_slv(opcode_type, 16#08#),
      883 => to_slv(opcode_type, 16#0F#),
      884 => to_slv(opcode_type, 16#0D#),
      885 => to_slv(opcode_type, 16#06#),
      886 => to_slv(opcode_type, 16#0A#),
      887 => to_slv(opcode_type, 16#0D#),
      888 => to_slv(opcode_type, 16#06#),
      889 => to_slv(opcode_type, 16#05#),
      890 => to_slv(opcode_type, 16#0D#),
      891 => to_slv(opcode_type, 16#01#),
      892 => to_slv(opcode_type, 16#0C#),
      893 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#07#),
      897 => to_slv(opcode_type, 16#06#),
      898 => to_slv(opcode_type, 16#06#),
      899 => to_slv(opcode_type, 16#02#),
      900 => to_slv(opcode_type, 16#11#),
      901 => to_slv(opcode_type, 16#04#),
      902 => to_slv(opcode_type, 16#0C#),
      903 => to_slv(opcode_type, 16#09#),
      904 => to_slv(opcode_type, 16#08#),
      905 => to_slv(opcode_type, 16#0E#),
      906 => to_slv(opcode_type, 16#0D#),
      907 => to_slv(opcode_type, 16#07#),
      908 => to_slv(opcode_type, 16#0C#),
      909 => to_slv(opcode_type, 16#47#),
      910 => to_slv(opcode_type, 16#06#),
      911 => to_slv(opcode_type, 16#09#),
      912 => to_slv(opcode_type, 16#09#),
      913 => to_slv(opcode_type, 16#0A#),
      914 => to_slv(opcode_type, 16#10#),
      915 => to_slv(opcode_type, 16#06#),
      916 => to_slv(opcode_type, 16#0D#),
      917 => to_slv(opcode_type, 16#0F#),
      918 => to_slv(opcode_type, 16#06#),
      919 => to_slv(opcode_type, 16#06#),
      920 => to_slv(opcode_type, 16#10#),
      921 => to_slv(opcode_type, 16#9B#),
      922 => to_slv(opcode_type, 16#09#),
      923 => to_slv(opcode_type, 16#0A#),
      924 => to_slv(opcode_type, 16#10#),
      925 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#09#),
      929 => to_slv(opcode_type, 16#06#),
      930 => to_slv(opcode_type, 16#09#),
      931 => to_slv(opcode_type, 16#01#),
      932 => to_slv(opcode_type, 16#0D#),
      933 => to_slv(opcode_type, 16#08#),
      934 => to_slv(opcode_type, 16#E7#),
      935 => to_slv(opcode_type, 16#0F#),
      936 => to_slv(opcode_type, 16#09#),
      937 => to_slv(opcode_type, 16#03#),
      938 => to_slv(opcode_type, 16#F9#),
      939 => to_slv(opcode_type, 16#07#),
      940 => to_slv(opcode_type, 16#0D#),
      941 => to_slv(opcode_type, 16#14#),
      942 => to_slv(opcode_type, 16#07#),
      943 => to_slv(opcode_type, 16#07#),
      944 => to_slv(opcode_type, 16#07#),
      945 => to_slv(opcode_type, 16#0B#),
      946 => to_slv(opcode_type, 16#10#),
      947 => to_slv(opcode_type, 16#08#),
      948 => to_slv(opcode_type, 16#0F#),
      949 => to_slv(opcode_type, 16#10#),
      950 => to_slv(opcode_type, 16#07#),
      951 => to_slv(opcode_type, 16#08#),
      952 => to_slv(opcode_type, 16#0C#),
      953 => to_slv(opcode_type, 16#EE#),
      954 => to_slv(opcode_type, 16#09#),
      955 => to_slv(opcode_type, 16#0D#),
      956 => to_slv(opcode_type, 16#0B#),
      957 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#08#),
      961 => to_slv(opcode_type, 16#08#),
      962 => to_slv(opcode_type, 16#06#),
      963 => to_slv(opcode_type, 16#09#),
      964 => to_slv(opcode_type, 16#5C#),
      965 => to_slv(opcode_type, 16#0F#),
      966 => to_slv(opcode_type, 16#07#),
      967 => to_slv(opcode_type, 16#0E#),
      968 => to_slv(opcode_type, 16#27#),
      969 => to_slv(opcode_type, 16#06#),
      970 => to_slv(opcode_type, 16#09#),
      971 => to_slv(opcode_type, 16#0D#),
      972 => to_slv(opcode_type, 16#11#),
      973 => to_slv(opcode_type, 16#05#),
      974 => to_slv(opcode_type, 16#11#),
      975 => to_slv(opcode_type, 16#06#),
      976 => to_slv(opcode_type, 16#08#),
      977 => to_slv(opcode_type, 16#06#),
      978 => to_slv(opcode_type, 16#0E#),
      979 => to_slv(opcode_type, 16#11#),
      980 => to_slv(opcode_type, 16#06#),
      981 => to_slv(opcode_type, 16#0D#),
      982 => to_slv(opcode_type, 16#0B#),
      983 => to_slv(opcode_type, 16#07#),
      984 => to_slv(opcode_type, 16#09#),
      985 => to_slv(opcode_type, 16#0F#),
      986 => to_slv(opcode_type, 16#10#),
      987 => to_slv(opcode_type, 16#05#),
      988 => to_slv(opcode_type, 16#10#),
      989 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#09#),
      993 => to_slv(opcode_type, 16#07#),
      994 => to_slv(opcode_type, 16#06#),
      995 => to_slv(opcode_type, 16#07#),
      996 => to_slv(opcode_type, 16#10#),
      997 => to_slv(opcode_type, 16#0B#),
      998 => to_slv(opcode_type, 16#09#),
      999 => to_slv(opcode_type, 16#0D#),
      1000 => to_slv(opcode_type, 16#0B#),
      1001 => to_slv(opcode_type, 16#08#),
      1002 => to_slv(opcode_type, 16#04#),
      1003 => to_slv(opcode_type, 16#11#),
      1004 => to_slv(opcode_type, 16#01#),
      1005 => to_slv(opcode_type, 16#0E#),
      1006 => to_slv(opcode_type, 16#07#),
      1007 => to_slv(opcode_type, 16#06#),
      1008 => to_slv(opcode_type, 16#07#),
      1009 => to_slv(opcode_type, 16#84#),
      1010 => to_slv(opcode_type, 16#31#),
      1011 => to_slv(opcode_type, 16#09#),
      1012 => to_slv(opcode_type, 16#0A#),
      1013 => to_slv(opcode_type, 16#0D#),
      1014 => to_slv(opcode_type, 16#06#),
      1015 => to_slv(opcode_type, 16#07#),
      1016 => to_slv(opcode_type, 16#0C#),
      1017 => to_slv(opcode_type, 16#13#),
      1018 => to_slv(opcode_type, 16#06#),
      1019 => to_slv(opcode_type, 16#0D#),
      1020 => to_slv(opcode_type, 16#0C#),
      1021 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#08#),
      1025 => to_slv(opcode_type, 16#07#),
      1026 => to_slv(opcode_type, 16#08#),
      1027 => to_slv(opcode_type, 16#04#),
      1028 => to_slv(opcode_type, 16#0D#),
      1029 => to_slv(opcode_type, 16#01#),
      1030 => to_slv(opcode_type, 16#0C#),
      1031 => to_slv(opcode_type, 16#09#),
      1032 => to_slv(opcode_type, 16#09#),
      1033 => to_slv(opcode_type, 16#0C#),
      1034 => to_slv(opcode_type, 16#11#),
      1035 => to_slv(opcode_type, 16#08#),
      1036 => to_slv(opcode_type, 16#10#),
      1037 => to_slv(opcode_type, 16#10#),
      1038 => to_slv(opcode_type, 16#07#),
      1039 => to_slv(opcode_type, 16#09#),
      1040 => to_slv(opcode_type, 16#09#),
      1041 => to_slv(opcode_type, 16#0D#),
      1042 => to_slv(opcode_type, 16#0C#),
      1043 => to_slv(opcode_type, 16#07#),
      1044 => to_slv(opcode_type, 16#0E#),
      1045 => to_slv(opcode_type, 16#8D#),
      1046 => to_slv(opcode_type, 16#08#),
      1047 => to_slv(opcode_type, 16#07#),
      1048 => to_slv(opcode_type, 16#0D#),
      1049 => to_slv(opcode_type, 16#0B#),
      1050 => to_slv(opcode_type, 16#09#),
      1051 => to_slv(opcode_type, 16#0E#),
      1052 => to_slv(opcode_type, 16#0E#),
      1053 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#07#),
      1057 => to_slv(opcode_type, 16#06#),
      1058 => to_slv(opcode_type, 16#08#),
      1059 => to_slv(opcode_type, 16#02#),
      1060 => to_slv(opcode_type, 16#11#),
      1061 => to_slv(opcode_type, 16#07#),
      1062 => to_slv(opcode_type, 16#EC#),
      1063 => to_slv(opcode_type, 16#3A#),
      1064 => to_slv(opcode_type, 16#06#),
      1065 => to_slv(opcode_type, 16#07#),
      1066 => to_slv(opcode_type, 16#0E#),
      1067 => to_slv(opcode_type, 16#0D#),
      1068 => to_slv(opcode_type, 16#08#),
      1069 => to_slv(opcode_type, 16#11#),
      1070 => to_slv(opcode_type, 16#AB#),
      1071 => to_slv(opcode_type, 16#07#),
      1072 => to_slv(opcode_type, 16#08#),
      1073 => to_slv(opcode_type, 16#03#),
      1074 => to_slv(opcode_type, 16#0A#),
      1075 => to_slv(opcode_type, 16#06#),
      1076 => to_slv(opcode_type, 16#0D#),
      1077 => to_slv(opcode_type, 16#0B#),
      1078 => to_slv(opcode_type, 16#09#),
      1079 => to_slv(opcode_type, 16#08#),
      1080 => to_slv(opcode_type, 16#0C#),
      1081 => to_slv(opcode_type, 16#0A#),
      1082 => to_slv(opcode_type, 16#06#),
      1083 => to_slv(opcode_type, 16#0F#),
      1084 => to_slv(opcode_type, 16#0E#),
      1085 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#09#),
      1089 => to_slv(opcode_type, 16#06#),
      1090 => to_slv(opcode_type, 16#08#),
      1091 => to_slv(opcode_type, 16#06#),
      1092 => to_slv(opcode_type, 16#0E#),
      1093 => to_slv(opcode_type, 16#0A#),
      1094 => to_slv(opcode_type, 16#05#),
      1095 => to_slv(opcode_type, 16#0A#),
      1096 => to_slv(opcode_type, 16#08#),
      1097 => to_slv(opcode_type, 16#01#),
      1098 => to_slv(opcode_type, 16#11#),
      1099 => to_slv(opcode_type, 16#08#),
      1100 => to_slv(opcode_type, 16#10#),
      1101 => to_slv(opcode_type, 16#0D#),
      1102 => to_slv(opcode_type, 16#06#),
      1103 => to_slv(opcode_type, 16#08#),
      1104 => to_slv(opcode_type, 16#07#),
      1105 => to_slv(opcode_type, 16#0B#),
      1106 => to_slv(opcode_type, 16#0E#),
      1107 => to_slv(opcode_type, 16#06#),
      1108 => to_slv(opcode_type, 16#10#),
      1109 => to_slv(opcode_type, 16#11#),
      1110 => to_slv(opcode_type, 16#09#),
      1111 => to_slv(opcode_type, 16#07#),
      1112 => to_slv(opcode_type, 16#10#),
      1113 => to_slv(opcode_type, 16#0A#),
      1114 => to_slv(opcode_type, 16#07#),
      1115 => to_slv(opcode_type, 16#0E#),
      1116 => to_slv(opcode_type, 16#56#),
      1117 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#09#),
      1121 => to_slv(opcode_type, 16#08#),
      1122 => to_slv(opcode_type, 16#08#),
      1123 => to_slv(opcode_type, 16#07#),
      1124 => to_slv(opcode_type, 16#0D#),
      1125 => to_slv(opcode_type, 16#97#),
      1126 => to_slv(opcode_type, 16#01#),
      1127 => to_slv(opcode_type, 16#0C#),
      1128 => to_slv(opcode_type, 16#09#),
      1129 => to_slv(opcode_type, 16#02#),
      1130 => to_slv(opcode_type, 16#0F#),
      1131 => to_slv(opcode_type, 16#06#),
      1132 => to_slv(opcode_type, 16#0C#),
      1133 => to_slv(opcode_type, 16#77#),
      1134 => to_slv(opcode_type, 16#09#),
      1135 => to_slv(opcode_type, 16#06#),
      1136 => to_slv(opcode_type, 16#08#),
      1137 => to_slv(opcode_type, 16#11#),
      1138 => to_slv(opcode_type, 16#0A#),
      1139 => to_slv(opcode_type, 16#07#),
      1140 => to_slv(opcode_type, 16#0E#),
      1141 => to_slv(opcode_type, 16#0B#),
      1142 => to_slv(opcode_type, 16#07#),
      1143 => to_slv(opcode_type, 16#09#),
      1144 => to_slv(opcode_type, 16#0E#),
      1145 => to_slv(opcode_type, 16#11#),
      1146 => to_slv(opcode_type, 16#08#),
      1147 => to_slv(opcode_type, 16#0C#),
      1148 => to_slv(opcode_type, 16#0E#),
      1149 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#08#),
      1153 => to_slv(opcode_type, 16#07#),
      1154 => to_slv(opcode_type, 16#09#),
      1155 => to_slv(opcode_type, 16#03#),
      1156 => to_slv(opcode_type, 16#0F#),
      1157 => to_slv(opcode_type, 16#08#),
      1158 => to_slv(opcode_type, 16#11#),
      1159 => to_slv(opcode_type, 16#11#),
      1160 => to_slv(opcode_type, 16#06#),
      1161 => to_slv(opcode_type, 16#02#),
      1162 => to_slv(opcode_type, 16#11#),
      1163 => to_slv(opcode_type, 16#09#),
      1164 => to_slv(opcode_type, 16#0B#),
      1165 => to_slv(opcode_type, 16#DB#),
      1166 => to_slv(opcode_type, 16#08#),
      1167 => to_slv(opcode_type, 16#06#),
      1168 => to_slv(opcode_type, 16#06#),
      1169 => to_slv(opcode_type, 16#0C#),
      1170 => to_slv(opcode_type, 16#10#),
      1171 => to_slv(opcode_type, 16#09#),
      1172 => to_slv(opcode_type, 16#0F#),
      1173 => to_slv(opcode_type, 16#10#),
      1174 => to_slv(opcode_type, 16#07#),
      1175 => to_slv(opcode_type, 16#09#),
      1176 => to_slv(opcode_type, 16#10#),
      1177 => to_slv(opcode_type, 16#0B#),
      1178 => to_slv(opcode_type, 16#07#),
      1179 => to_slv(opcode_type, 16#0A#),
      1180 => to_slv(opcode_type, 16#0F#),
      1181 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#07#),
      1185 => to_slv(opcode_type, 16#07#),
      1186 => to_slv(opcode_type, 16#09#),
      1187 => to_slv(opcode_type, 16#06#),
      1188 => to_slv(opcode_type, 16#67#),
      1189 => to_slv(opcode_type, 16#0D#),
      1190 => to_slv(opcode_type, 16#02#),
      1191 => to_slv(opcode_type, 16#11#),
      1192 => to_slv(opcode_type, 16#08#),
      1193 => to_slv(opcode_type, 16#01#),
      1194 => to_slv(opcode_type, 16#11#),
      1195 => to_slv(opcode_type, 16#08#),
      1196 => to_slv(opcode_type, 16#0F#),
      1197 => to_slv(opcode_type, 16#0D#),
      1198 => to_slv(opcode_type, 16#08#),
      1199 => to_slv(opcode_type, 16#07#),
      1200 => to_slv(opcode_type, 16#08#),
      1201 => to_slv(opcode_type, 16#0D#),
      1202 => to_slv(opcode_type, 16#0C#),
      1203 => to_slv(opcode_type, 16#06#),
      1204 => to_slv(opcode_type, 16#0F#),
      1205 => to_slv(opcode_type, 16#10#),
      1206 => to_slv(opcode_type, 16#09#),
      1207 => to_slv(opcode_type, 16#06#),
      1208 => to_slv(opcode_type, 16#0F#),
      1209 => to_slv(opcode_type, 16#0C#),
      1210 => to_slv(opcode_type, 16#07#),
      1211 => to_slv(opcode_type, 16#0A#),
      1212 => to_slv(opcode_type, 16#0B#),
      1213 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#08#),
      1217 => to_slv(opcode_type, 16#06#),
      1218 => to_slv(opcode_type, 16#08#),
      1219 => to_slv(opcode_type, 16#05#),
      1220 => to_slv(opcode_type, 16#0E#),
      1221 => to_slv(opcode_type, 16#09#),
      1222 => to_slv(opcode_type, 16#FE#),
      1223 => to_slv(opcode_type, 16#96#),
      1224 => to_slv(opcode_type, 16#08#),
      1225 => to_slv(opcode_type, 16#09#),
      1226 => to_slv(opcode_type, 16#0F#),
      1227 => to_slv(opcode_type, 16#0D#),
      1228 => to_slv(opcode_type, 16#05#),
      1229 => to_slv(opcode_type, 16#11#),
      1230 => to_slv(opcode_type, 16#09#),
      1231 => to_slv(opcode_type, 16#07#),
      1232 => to_slv(opcode_type, 16#09#),
      1233 => to_slv(opcode_type, 16#11#),
      1234 => to_slv(opcode_type, 16#0C#),
      1235 => to_slv(opcode_type, 16#07#),
      1236 => to_slv(opcode_type, 16#89#),
      1237 => to_slv(opcode_type, 16#0C#),
      1238 => to_slv(opcode_type, 16#07#),
      1239 => to_slv(opcode_type, 16#08#),
      1240 => to_slv(opcode_type, 16#0C#),
      1241 => to_slv(opcode_type, 16#10#),
      1242 => to_slv(opcode_type, 16#09#),
      1243 => to_slv(opcode_type, 16#0E#),
      1244 => to_slv(opcode_type, 16#10#),
      1245 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#06#),
      1249 => to_slv(opcode_type, 16#08#),
      1250 => to_slv(opcode_type, 16#07#),
      1251 => to_slv(opcode_type, 16#02#),
      1252 => to_slv(opcode_type, 16#0A#),
      1253 => to_slv(opcode_type, 16#02#),
      1254 => to_slv(opcode_type, 16#0F#),
      1255 => to_slv(opcode_type, 16#07#),
      1256 => to_slv(opcode_type, 16#07#),
      1257 => to_slv(opcode_type, 16#0B#),
      1258 => to_slv(opcode_type, 16#0B#),
      1259 => to_slv(opcode_type, 16#07#),
      1260 => to_slv(opcode_type, 16#0F#),
      1261 => to_slv(opcode_type, 16#0C#),
      1262 => to_slv(opcode_type, 16#07#),
      1263 => to_slv(opcode_type, 16#08#),
      1264 => to_slv(opcode_type, 16#07#),
      1265 => to_slv(opcode_type, 16#0E#),
      1266 => to_slv(opcode_type, 16#0D#),
      1267 => to_slv(opcode_type, 16#06#),
      1268 => to_slv(opcode_type, 16#BD#),
      1269 => to_slv(opcode_type, 16#1D#),
      1270 => to_slv(opcode_type, 16#07#),
      1271 => to_slv(opcode_type, 16#07#),
      1272 => to_slv(opcode_type, 16#0C#),
      1273 => to_slv(opcode_type, 16#0E#),
      1274 => to_slv(opcode_type, 16#09#),
      1275 => to_slv(opcode_type, 16#0A#),
      1276 => to_slv(opcode_type, 16#0F#),
      1277 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#09#),
      1281 => to_slv(opcode_type, 16#09#),
      1282 => to_slv(opcode_type, 16#09#),
      1283 => to_slv(opcode_type, 16#02#),
      1284 => to_slv(opcode_type, 16#10#),
      1285 => to_slv(opcode_type, 16#04#),
      1286 => to_slv(opcode_type, 16#0D#),
      1287 => to_slv(opcode_type, 16#08#),
      1288 => to_slv(opcode_type, 16#08#),
      1289 => to_slv(opcode_type, 16#0A#),
      1290 => to_slv(opcode_type, 16#C6#),
      1291 => to_slv(opcode_type, 16#08#),
      1292 => to_slv(opcode_type, 16#0D#),
      1293 => to_slv(opcode_type, 16#0C#),
      1294 => to_slv(opcode_type, 16#08#),
      1295 => to_slv(opcode_type, 16#07#),
      1296 => to_slv(opcode_type, 16#07#),
      1297 => to_slv(opcode_type, 16#0E#),
      1298 => to_slv(opcode_type, 16#0C#),
      1299 => to_slv(opcode_type, 16#07#),
      1300 => to_slv(opcode_type, 16#0D#),
      1301 => to_slv(opcode_type, 16#0C#),
      1302 => to_slv(opcode_type, 16#09#),
      1303 => to_slv(opcode_type, 16#08#),
      1304 => to_slv(opcode_type, 16#0F#),
      1305 => to_slv(opcode_type, 16#11#),
      1306 => to_slv(opcode_type, 16#07#),
      1307 => to_slv(opcode_type, 16#0A#),
      1308 => to_slv(opcode_type, 16#70#),
      1309 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#08#),
      1313 => to_slv(opcode_type, 16#09#),
      1314 => to_slv(opcode_type, 16#06#),
      1315 => to_slv(opcode_type, 16#01#),
      1316 => to_slv(opcode_type, 16#0F#),
      1317 => to_slv(opcode_type, 16#04#),
      1318 => to_slv(opcode_type, 16#0E#),
      1319 => to_slv(opcode_type, 16#07#),
      1320 => to_slv(opcode_type, 16#07#),
      1321 => to_slv(opcode_type, 16#11#),
      1322 => to_slv(opcode_type, 16#54#),
      1323 => to_slv(opcode_type, 16#08#),
      1324 => to_slv(opcode_type, 16#10#),
      1325 => to_slv(opcode_type, 16#0E#),
      1326 => to_slv(opcode_type, 16#08#),
      1327 => to_slv(opcode_type, 16#06#),
      1328 => to_slv(opcode_type, 16#09#),
      1329 => to_slv(opcode_type, 16#0D#),
      1330 => to_slv(opcode_type, 16#0E#),
      1331 => to_slv(opcode_type, 16#07#),
      1332 => to_slv(opcode_type, 16#0C#),
      1333 => to_slv(opcode_type, 16#11#),
      1334 => to_slv(opcode_type, 16#07#),
      1335 => to_slv(opcode_type, 16#07#),
      1336 => to_slv(opcode_type, 16#11#),
      1337 => to_slv(opcode_type, 16#10#),
      1338 => to_slv(opcode_type, 16#08#),
      1339 => to_slv(opcode_type, 16#0B#),
      1340 => to_slv(opcode_type, 16#10#),
      1341 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#07#),
      1345 => to_slv(opcode_type, 16#07#),
      1346 => to_slv(opcode_type, 16#08#),
      1347 => to_slv(opcode_type, 16#02#),
      1348 => to_slv(opcode_type, 16#0F#),
      1349 => to_slv(opcode_type, 16#06#),
      1350 => to_slv(opcode_type, 16#0C#),
      1351 => to_slv(opcode_type, 16#0A#),
      1352 => to_slv(opcode_type, 16#06#),
      1353 => to_slv(opcode_type, 16#07#),
      1354 => to_slv(opcode_type, 16#0C#),
      1355 => to_slv(opcode_type, 16#0B#),
      1356 => to_slv(opcode_type, 16#09#),
      1357 => to_slv(opcode_type, 16#0E#),
      1358 => to_slv(opcode_type, 16#10#),
      1359 => to_slv(opcode_type, 16#08#),
      1360 => to_slv(opcode_type, 16#07#),
      1361 => to_slv(opcode_type, 16#01#),
      1362 => to_slv(opcode_type, 16#0D#),
      1363 => to_slv(opcode_type, 16#06#),
      1364 => to_slv(opcode_type, 16#0E#),
      1365 => to_slv(opcode_type, 16#10#),
      1366 => to_slv(opcode_type, 16#08#),
      1367 => to_slv(opcode_type, 16#06#),
      1368 => to_slv(opcode_type, 16#0D#),
      1369 => to_slv(opcode_type, 16#0C#),
      1370 => to_slv(opcode_type, 16#06#),
      1371 => to_slv(opcode_type, 16#0C#),
      1372 => to_slv(opcode_type, 16#0A#),
      1373 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#07#),
      1377 => to_slv(opcode_type, 16#06#),
      1378 => to_slv(opcode_type, 16#08#),
      1379 => to_slv(opcode_type, 16#02#),
      1380 => to_slv(opcode_type, 16#0D#),
      1381 => to_slv(opcode_type, 16#09#),
      1382 => to_slv(opcode_type, 16#0A#),
      1383 => to_slv(opcode_type, 16#11#),
      1384 => to_slv(opcode_type, 16#06#),
      1385 => to_slv(opcode_type, 16#09#),
      1386 => to_slv(opcode_type, 16#0E#),
      1387 => to_slv(opcode_type, 16#10#),
      1388 => to_slv(opcode_type, 16#02#),
      1389 => to_slv(opcode_type, 16#0A#),
      1390 => to_slv(opcode_type, 16#07#),
      1391 => to_slv(opcode_type, 16#06#),
      1392 => to_slv(opcode_type, 16#06#),
      1393 => to_slv(opcode_type, 16#0B#),
      1394 => to_slv(opcode_type, 16#30#),
      1395 => to_slv(opcode_type, 16#06#),
      1396 => to_slv(opcode_type, 16#0F#),
      1397 => to_slv(opcode_type, 16#0F#),
      1398 => to_slv(opcode_type, 16#09#),
      1399 => to_slv(opcode_type, 16#07#),
      1400 => to_slv(opcode_type, 16#0C#),
      1401 => to_slv(opcode_type, 16#10#),
      1402 => to_slv(opcode_type, 16#06#),
      1403 => to_slv(opcode_type, 16#4C#),
      1404 => to_slv(opcode_type, 16#10#),
      1405 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#08#),
      1409 => to_slv(opcode_type, 16#07#),
      1410 => to_slv(opcode_type, 16#08#),
      1411 => to_slv(opcode_type, 16#07#),
      1412 => to_slv(opcode_type, 16#0B#),
      1413 => to_slv(opcode_type, 16#0E#),
      1414 => to_slv(opcode_type, 16#09#),
      1415 => to_slv(opcode_type, 16#0C#),
      1416 => to_slv(opcode_type, 16#0B#),
      1417 => to_slv(opcode_type, 16#07#),
      1418 => to_slv(opcode_type, 16#09#),
      1419 => to_slv(opcode_type, 16#CA#),
      1420 => to_slv(opcode_type, 16#73#),
      1421 => to_slv(opcode_type, 16#08#),
      1422 => to_slv(opcode_type, 16#0B#),
      1423 => to_slv(opcode_type, 16#0B#),
      1424 => to_slv(opcode_type, 16#09#),
      1425 => to_slv(opcode_type, 16#08#),
      1426 => to_slv(opcode_type, 16#08#),
      1427 => to_slv(opcode_type, 16#0B#),
      1428 => to_slv(opcode_type, 16#0C#),
      1429 => to_slv(opcode_type, 16#05#),
      1430 => to_slv(opcode_type, 16#0C#),
      1431 => to_slv(opcode_type, 16#06#),
      1432 => to_slv(opcode_type, 16#08#),
      1433 => to_slv(opcode_type, 16#0C#),
      1434 => to_slv(opcode_type, 16#10#),
      1435 => to_slv(opcode_type, 16#01#),
      1436 => to_slv(opcode_type, 16#0B#),
      1437 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#06#),
      1441 => to_slv(opcode_type, 16#07#),
      1442 => to_slv(opcode_type, 16#08#),
      1443 => to_slv(opcode_type, 16#09#),
      1444 => to_slv(opcode_type, 16#0B#),
      1445 => to_slv(opcode_type, 16#0E#),
      1446 => to_slv(opcode_type, 16#08#),
      1447 => to_slv(opcode_type, 16#0F#),
      1448 => to_slv(opcode_type, 16#0C#),
      1449 => to_slv(opcode_type, 16#08#),
      1450 => to_slv(opcode_type, 16#03#),
      1451 => to_slv(opcode_type, 16#11#),
      1452 => to_slv(opcode_type, 16#02#),
      1453 => to_slv(opcode_type, 16#0A#),
      1454 => to_slv(opcode_type, 16#09#),
      1455 => to_slv(opcode_type, 16#08#),
      1456 => to_slv(opcode_type, 16#06#),
      1457 => to_slv(opcode_type, 16#10#),
      1458 => to_slv(opcode_type, 16#0F#),
      1459 => to_slv(opcode_type, 16#08#),
      1460 => to_slv(opcode_type, 16#0F#),
      1461 => to_slv(opcode_type, 16#11#),
      1462 => to_slv(opcode_type, 16#09#),
      1463 => to_slv(opcode_type, 16#09#),
      1464 => to_slv(opcode_type, 16#0B#),
      1465 => to_slv(opcode_type, 16#11#),
      1466 => to_slv(opcode_type, 16#09#),
      1467 => to_slv(opcode_type, 16#0A#),
      1468 => to_slv(opcode_type, 16#0F#),
      1469 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#06#),
      1473 => to_slv(opcode_type, 16#06#),
      1474 => to_slv(opcode_type, 16#09#),
      1475 => to_slv(opcode_type, 16#01#),
      1476 => to_slv(opcode_type, 16#3F#),
      1477 => to_slv(opcode_type, 16#09#),
      1478 => to_slv(opcode_type, 16#0E#),
      1479 => to_slv(opcode_type, 16#0D#),
      1480 => to_slv(opcode_type, 16#08#),
      1481 => to_slv(opcode_type, 16#07#),
      1482 => to_slv(opcode_type, 16#0E#),
      1483 => to_slv(opcode_type, 16#0C#),
      1484 => to_slv(opcode_type, 16#09#),
      1485 => to_slv(opcode_type, 16#0C#),
      1486 => to_slv(opcode_type, 16#0D#),
      1487 => to_slv(opcode_type, 16#09#),
      1488 => to_slv(opcode_type, 16#06#),
      1489 => to_slv(opcode_type, 16#05#),
      1490 => to_slv(opcode_type, 16#0C#),
      1491 => to_slv(opcode_type, 16#06#),
      1492 => to_slv(opcode_type, 16#0F#),
      1493 => to_slv(opcode_type, 16#0E#),
      1494 => to_slv(opcode_type, 16#06#),
      1495 => to_slv(opcode_type, 16#09#),
      1496 => to_slv(opcode_type, 16#0E#),
      1497 => to_slv(opcode_type, 16#0E#),
      1498 => to_slv(opcode_type, 16#07#),
      1499 => to_slv(opcode_type, 16#0D#),
      1500 => to_slv(opcode_type, 16#0C#),
      1501 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#07#),
      1505 => to_slv(opcode_type, 16#06#),
      1506 => to_slv(opcode_type, 16#06#),
      1507 => to_slv(opcode_type, 16#08#),
      1508 => to_slv(opcode_type, 16#28#),
      1509 => to_slv(opcode_type, 16#5B#),
      1510 => to_slv(opcode_type, 16#08#),
      1511 => to_slv(opcode_type, 16#0E#),
      1512 => to_slv(opcode_type, 16#0E#),
      1513 => to_slv(opcode_type, 16#07#),
      1514 => to_slv(opcode_type, 16#01#),
      1515 => to_slv(opcode_type, 16#0D#),
      1516 => to_slv(opcode_type, 16#03#),
      1517 => to_slv(opcode_type, 16#11#),
      1518 => to_slv(opcode_type, 16#07#),
      1519 => to_slv(opcode_type, 16#06#),
      1520 => to_slv(opcode_type, 16#08#),
      1521 => to_slv(opcode_type, 16#0A#),
      1522 => to_slv(opcode_type, 16#24#),
      1523 => to_slv(opcode_type, 16#08#),
      1524 => to_slv(opcode_type, 16#10#),
      1525 => to_slv(opcode_type, 16#0E#),
      1526 => to_slv(opcode_type, 16#09#),
      1527 => to_slv(opcode_type, 16#08#),
      1528 => to_slv(opcode_type, 16#11#),
      1529 => to_slv(opcode_type, 16#51#),
      1530 => to_slv(opcode_type, 16#09#),
      1531 => to_slv(opcode_type, 16#11#),
      1532 => to_slv(opcode_type, 16#0D#),
      1533 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#07#),
      1537 => to_slv(opcode_type, 16#07#),
      1538 => to_slv(opcode_type, 16#08#),
      1539 => to_slv(opcode_type, 16#02#),
      1540 => to_slv(opcode_type, 16#0B#),
      1541 => to_slv(opcode_type, 16#06#),
      1542 => to_slv(opcode_type, 16#82#),
      1543 => to_slv(opcode_type, 16#0B#),
      1544 => to_slv(opcode_type, 16#08#),
      1545 => to_slv(opcode_type, 16#02#),
      1546 => to_slv(opcode_type, 16#0B#),
      1547 => to_slv(opcode_type, 16#07#),
      1548 => to_slv(opcode_type, 16#0E#),
      1549 => to_slv(opcode_type, 16#0C#),
      1550 => to_slv(opcode_type, 16#07#),
      1551 => to_slv(opcode_type, 16#08#),
      1552 => to_slv(opcode_type, 16#08#),
      1553 => to_slv(opcode_type, 16#11#),
      1554 => to_slv(opcode_type, 16#5E#),
      1555 => to_slv(opcode_type, 16#06#),
      1556 => to_slv(opcode_type, 16#0C#),
      1557 => to_slv(opcode_type, 16#8A#),
      1558 => to_slv(opcode_type, 16#08#),
      1559 => to_slv(opcode_type, 16#09#),
      1560 => to_slv(opcode_type, 16#10#),
      1561 => to_slv(opcode_type, 16#0D#),
      1562 => to_slv(opcode_type, 16#09#),
      1563 => to_slv(opcode_type, 16#0F#),
      1564 => to_slv(opcode_type, 16#10#),
      1565 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#08#),
      1569 => to_slv(opcode_type, 16#06#),
      1570 => to_slv(opcode_type, 16#06#),
      1571 => to_slv(opcode_type, 16#03#),
      1572 => to_slv(opcode_type, 16#11#),
      1573 => to_slv(opcode_type, 16#01#),
      1574 => to_slv(opcode_type, 16#0F#),
      1575 => to_slv(opcode_type, 16#07#),
      1576 => to_slv(opcode_type, 16#06#),
      1577 => to_slv(opcode_type, 16#0D#),
      1578 => to_slv(opcode_type, 16#0F#),
      1579 => to_slv(opcode_type, 16#07#),
      1580 => to_slv(opcode_type, 16#2F#),
      1581 => to_slv(opcode_type, 16#0E#),
      1582 => to_slv(opcode_type, 16#09#),
      1583 => to_slv(opcode_type, 16#08#),
      1584 => to_slv(opcode_type, 16#08#),
      1585 => to_slv(opcode_type, 16#0A#),
      1586 => to_slv(opcode_type, 16#10#),
      1587 => to_slv(opcode_type, 16#09#),
      1588 => to_slv(opcode_type, 16#0C#),
      1589 => to_slv(opcode_type, 16#0D#),
      1590 => to_slv(opcode_type, 16#09#),
      1591 => to_slv(opcode_type, 16#07#),
      1592 => to_slv(opcode_type, 16#0F#),
      1593 => to_slv(opcode_type, 16#10#),
      1594 => to_slv(opcode_type, 16#08#),
      1595 => to_slv(opcode_type, 16#0E#),
      1596 => to_slv(opcode_type, 16#0A#),
      1597 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#08#),
      1602 => to_slv(opcode_type, 16#08#),
      1603 => to_slv(opcode_type, 16#04#),
      1604 => to_slv(opcode_type, 16#0E#),
      1605 => to_slv(opcode_type, 16#05#),
      1606 => to_slv(opcode_type, 16#0E#),
      1607 => to_slv(opcode_type, 16#07#),
      1608 => to_slv(opcode_type, 16#07#),
      1609 => to_slv(opcode_type, 16#5C#),
      1610 => to_slv(opcode_type, 16#11#),
      1611 => to_slv(opcode_type, 16#09#),
      1612 => to_slv(opcode_type, 16#10#),
      1613 => to_slv(opcode_type, 16#FF#),
      1614 => to_slv(opcode_type, 16#08#),
      1615 => to_slv(opcode_type, 16#07#),
      1616 => to_slv(opcode_type, 16#07#),
      1617 => to_slv(opcode_type, 16#0C#),
      1618 => to_slv(opcode_type, 16#0C#),
      1619 => to_slv(opcode_type, 16#09#),
      1620 => to_slv(opcode_type, 16#0C#),
      1621 => to_slv(opcode_type, 16#0B#),
      1622 => to_slv(opcode_type, 16#08#),
      1623 => to_slv(opcode_type, 16#08#),
      1624 => to_slv(opcode_type, 16#0C#),
      1625 => to_slv(opcode_type, 16#87#),
      1626 => to_slv(opcode_type, 16#07#),
      1627 => to_slv(opcode_type, 16#0C#),
      1628 => to_slv(opcode_type, 16#0C#),
      1629 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#08#),
      1633 => to_slv(opcode_type, 16#07#),
      1634 => to_slv(opcode_type, 16#06#),
      1635 => to_slv(opcode_type, 16#04#),
      1636 => to_slv(opcode_type, 16#0F#),
      1637 => to_slv(opcode_type, 16#09#),
      1638 => to_slv(opcode_type, 16#0D#),
      1639 => to_slv(opcode_type, 16#0F#),
      1640 => to_slv(opcode_type, 16#06#),
      1641 => to_slv(opcode_type, 16#08#),
      1642 => to_slv(opcode_type, 16#10#),
      1643 => to_slv(opcode_type, 16#C1#),
      1644 => to_slv(opcode_type, 16#04#),
      1645 => to_slv(opcode_type, 16#0F#),
      1646 => to_slv(opcode_type, 16#07#),
      1647 => to_slv(opcode_type, 16#09#),
      1648 => to_slv(opcode_type, 16#07#),
      1649 => to_slv(opcode_type, 16#11#),
      1650 => to_slv(opcode_type, 16#39#),
      1651 => to_slv(opcode_type, 16#08#),
      1652 => to_slv(opcode_type, 16#0A#),
      1653 => to_slv(opcode_type, 16#11#),
      1654 => to_slv(opcode_type, 16#09#),
      1655 => to_slv(opcode_type, 16#09#),
      1656 => to_slv(opcode_type, 16#10#),
      1657 => to_slv(opcode_type, 16#11#),
      1658 => to_slv(opcode_type, 16#08#),
      1659 => to_slv(opcode_type, 16#0C#),
      1660 => to_slv(opcode_type, 16#0F#),
      1661 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#08#),
      1665 => to_slv(opcode_type, 16#09#),
      1666 => to_slv(opcode_type, 16#09#),
      1667 => to_slv(opcode_type, 16#05#),
      1668 => to_slv(opcode_type, 16#10#),
      1669 => to_slv(opcode_type, 16#01#),
      1670 => to_slv(opcode_type, 16#1E#),
      1671 => to_slv(opcode_type, 16#06#),
      1672 => to_slv(opcode_type, 16#08#),
      1673 => to_slv(opcode_type, 16#0E#),
      1674 => to_slv(opcode_type, 16#0E#),
      1675 => to_slv(opcode_type, 16#06#),
      1676 => to_slv(opcode_type, 16#0B#),
      1677 => to_slv(opcode_type, 16#0F#),
      1678 => to_slv(opcode_type, 16#06#),
      1679 => to_slv(opcode_type, 16#06#),
      1680 => to_slv(opcode_type, 16#09#),
      1681 => to_slv(opcode_type, 16#0A#),
      1682 => to_slv(opcode_type, 16#0C#),
      1683 => to_slv(opcode_type, 16#07#),
      1684 => to_slv(opcode_type, 16#10#),
      1685 => to_slv(opcode_type, 16#8E#),
      1686 => to_slv(opcode_type, 16#09#),
      1687 => to_slv(opcode_type, 16#09#),
      1688 => to_slv(opcode_type, 16#0F#),
      1689 => to_slv(opcode_type, 16#AB#),
      1690 => to_slv(opcode_type, 16#07#),
      1691 => to_slv(opcode_type, 16#0E#),
      1692 => to_slv(opcode_type, 16#10#),
      1693 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#06#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#07#),
      1699 => to_slv(opcode_type, 16#02#),
      1700 => to_slv(opcode_type, 16#C7#),
      1701 => to_slv(opcode_type, 16#06#),
      1702 => to_slv(opcode_type, 16#0E#),
      1703 => to_slv(opcode_type, 16#0A#),
      1704 => to_slv(opcode_type, 16#07#),
      1705 => to_slv(opcode_type, 16#05#),
      1706 => to_slv(opcode_type, 16#0A#),
      1707 => to_slv(opcode_type, 16#07#),
      1708 => to_slv(opcode_type, 16#10#),
      1709 => to_slv(opcode_type, 16#0C#),
      1710 => to_slv(opcode_type, 16#06#),
      1711 => to_slv(opcode_type, 16#09#),
      1712 => to_slv(opcode_type, 16#06#),
      1713 => to_slv(opcode_type, 16#0E#),
      1714 => to_slv(opcode_type, 16#76#),
      1715 => to_slv(opcode_type, 16#07#),
      1716 => to_slv(opcode_type, 16#10#),
      1717 => to_slv(opcode_type, 16#10#),
      1718 => to_slv(opcode_type, 16#09#),
      1719 => to_slv(opcode_type, 16#09#),
      1720 => to_slv(opcode_type, 16#0B#),
      1721 => to_slv(opcode_type, 16#10#),
      1722 => to_slv(opcode_type, 16#07#),
      1723 => to_slv(opcode_type, 16#11#),
      1724 => to_slv(opcode_type, 16#0A#),
      1725 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#07#),
      1729 => to_slv(opcode_type, 16#06#),
      1730 => to_slv(opcode_type, 16#07#),
      1731 => to_slv(opcode_type, 16#03#),
      1732 => to_slv(opcode_type, 16#0C#),
      1733 => to_slv(opcode_type, 16#08#),
      1734 => to_slv(opcode_type, 16#0B#),
      1735 => to_slv(opcode_type, 16#10#),
      1736 => to_slv(opcode_type, 16#09#),
      1737 => to_slv(opcode_type, 16#07#),
      1738 => to_slv(opcode_type, 16#0D#),
      1739 => to_slv(opcode_type, 16#0E#),
      1740 => to_slv(opcode_type, 16#02#),
      1741 => to_slv(opcode_type, 16#11#),
      1742 => to_slv(opcode_type, 16#07#),
      1743 => to_slv(opcode_type, 16#09#),
      1744 => to_slv(opcode_type, 16#06#),
      1745 => to_slv(opcode_type, 16#0E#),
      1746 => to_slv(opcode_type, 16#A3#),
      1747 => to_slv(opcode_type, 16#08#),
      1748 => to_slv(opcode_type, 16#10#),
      1749 => to_slv(opcode_type, 16#0C#),
      1750 => to_slv(opcode_type, 16#06#),
      1751 => to_slv(opcode_type, 16#06#),
      1752 => to_slv(opcode_type, 16#0D#),
      1753 => to_slv(opcode_type, 16#10#),
      1754 => to_slv(opcode_type, 16#06#),
      1755 => to_slv(opcode_type, 16#0C#),
      1756 => to_slv(opcode_type, 16#92#),
      1757 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#08#),
      1761 => to_slv(opcode_type, 16#09#),
      1762 => to_slv(opcode_type, 16#09#),
      1763 => to_slv(opcode_type, 16#04#),
      1764 => to_slv(opcode_type, 16#28#),
      1765 => to_slv(opcode_type, 16#03#),
      1766 => to_slv(opcode_type, 16#0E#),
      1767 => to_slv(opcode_type, 16#07#),
      1768 => to_slv(opcode_type, 16#06#),
      1769 => to_slv(opcode_type, 16#10#),
      1770 => to_slv(opcode_type, 16#11#),
      1771 => to_slv(opcode_type, 16#08#),
      1772 => to_slv(opcode_type, 16#10#),
      1773 => to_slv(opcode_type, 16#0C#),
      1774 => to_slv(opcode_type, 16#06#),
      1775 => to_slv(opcode_type, 16#09#),
      1776 => to_slv(opcode_type, 16#09#),
      1777 => to_slv(opcode_type, 16#7D#),
      1778 => to_slv(opcode_type, 16#0C#),
      1779 => to_slv(opcode_type, 16#09#),
      1780 => to_slv(opcode_type, 16#10#),
      1781 => to_slv(opcode_type, 16#EC#),
      1782 => to_slv(opcode_type, 16#09#),
      1783 => to_slv(opcode_type, 16#09#),
      1784 => to_slv(opcode_type, 16#0A#),
      1785 => to_slv(opcode_type, 16#0A#),
      1786 => to_slv(opcode_type, 16#07#),
      1787 => to_slv(opcode_type, 16#11#),
      1788 => to_slv(opcode_type, 16#0C#),
      1789 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#08#),
      1793 => to_slv(opcode_type, 16#06#),
      1794 => to_slv(opcode_type, 16#08#),
      1795 => to_slv(opcode_type, 16#02#),
      1796 => to_slv(opcode_type, 16#0E#),
      1797 => to_slv(opcode_type, 16#01#),
      1798 => to_slv(opcode_type, 16#0E#),
      1799 => to_slv(opcode_type, 16#06#),
      1800 => to_slv(opcode_type, 16#08#),
      1801 => to_slv(opcode_type, 16#0B#),
      1802 => to_slv(opcode_type, 16#0D#),
      1803 => to_slv(opcode_type, 16#07#),
      1804 => to_slv(opcode_type, 16#0C#),
      1805 => to_slv(opcode_type, 16#0B#),
      1806 => to_slv(opcode_type, 16#08#),
      1807 => to_slv(opcode_type, 16#09#),
      1808 => to_slv(opcode_type, 16#09#),
      1809 => to_slv(opcode_type, 16#0B#),
      1810 => to_slv(opcode_type, 16#11#),
      1811 => to_slv(opcode_type, 16#09#),
      1812 => to_slv(opcode_type, 16#86#),
      1813 => to_slv(opcode_type, 16#0C#),
      1814 => to_slv(opcode_type, 16#06#),
      1815 => to_slv(opcode_type, 16#06#),
      1816 => to_slv(opcode_type, 16#0E#),
      1817 => to_slv(opcode_type, 16#0A#),
      1818 => to_slv(opcode_type, 16#09#),
      1819 => to_slv(opcode_type, 16#0E#),
      1820 => to_slv(opcode_type, 16#0E#),
      1821 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#08#),
      1825 => to_slv(opcode_type, 16#09#),
      1826 => to_slv(opcode_type, 16#06#),
      1827 => to_slv(opcode_type, 16#05#),
      1828 => to_slv(opcode_type, 16#0A#),
      1829 => to_slv(opcode_type, 16#06#),
      1830 => to_slv(opcode_type, 16#AA#),
      1831 => to_slv(opcode_type, 16#0D#),
      1832 => to_slv(opcode_type, 16#06#),
      1833 => to_slv(opcode_type, 16#01#),
      1834 => to_slv(opcode_type, 16#11#),
      1835 => to_slv(opcode_type, 16#08#),
      1836 => to_slv(opcode_type, 16#B7#),
      1837 => to_slv(opcode_type, 16#0F#),
      1838 => to_slv(opcode_type, 16#07#),
      1839 => to_slv(opcode_type, 16#08#),
      1840 => to_slv(opcode_type, 16#09#),
      1841 => to_slv(opcode_type, 16#0B#),
      1842 => to_slv(opcode_type, 16#BB#),
      1843 => to_slv(opcode_type, 16#07#),
      1844 => to_slv(opcode_type, 16#10#),
      1845 => to_slv(opcode_type, 16#0F#),
      1846 => to_slv(opcode_type, 16#07#),
      1847 => to_slv(opcode_type, 16#06#),
      1848 => to_slv(opcode_type, 16#0A#),
      1849 => to_slv(opcode_type, 16#0F#),
      1850 => to_slv(opcode_type, 16#09#),
      1851 => to_slv(opcode_type, 16#0C#),
      1852 => to_slv(opcode_type, 16#0C#),
      1853 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#08#),
      1857 => to_slv(opcode_type, 16#08#),
      1858 => to_slv(opcode_type, 16#06#),
      1859 => to_slv(opcode_type, 16#06#),
      1860 => to_slv(opcode_type, 16#0D#),
      1861 => to_slv(opcode_type, 16#0F#),
      1862 => to_slv(opcode_type, 16#07#),
      1863 => to_slv(opcode_type, 16#0B#),
      1864 => to_slv(opcode_type, 16#0F#),
      1865 => to_slv(opcode_type, 16#06#),
      1866 => to_slv(opcode_type, 16#01#),
      1867 => to_slv(opcode_type, 16#0F#),
      1868 => to_slv(opcode_type, 16#01#),
      1869 => to_slv(opcode_type, 16#0E#),
      1870 => to_slv(opcode_type, 16#07#),
      1871 => to_slv(opcode_type, 16#06#),
      1872 => to_slv(opcode_type, 16#07#),
      1873 => to_slv(opcode_type, 16#0B#),
      1874 => to_slv(opcode_type, 16#0E#),
      1875 => to_slv(opcode_type, 16#09#),
      1876 => to_slv(opcode_type, 16#0F#),
      1877 => to_slv(opcode_type, 16#0D#),
      1878 => to_slv(opcode_type, 16#09#),
      1879 => to_slv(opcode_type, 16#07#),
      1880 => to_slv(opcode_type, 16#0F#),
      1881 => to_slv(opcode_type, 16#0A#),
      1882 => to_slv(opcode_type, 16#06#),
      1883 => to_slv(opcode_type, 16#10#),
      1884 => to_slv(opcode_type, 16#E1#),
      1885 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#09#),
      1889 => to_slv(opcode_type, 16#08#),
      1890 => to_slv(opcode_type, 16#09#),
      1891 => to_slv(opcode_type, 16#08#),
      1892 => to_slv(opcode_type, 16#0B#),
      1893 => to_slv(opcode_type, 16#0D#),
      1894 => to_slv(opcode_type, 16#01#),
      1895 => to_slv(opcode_type, 16#0C#),
      1896 => to_slv(opcode_type, 16#08#),
      1897 => to_slv(opcode_type, 16#06#),
      1898 => to_slv(opcode_type, 16#0A#),
      1899 => to_slv(opcode_type, 16#10#),
      1900 => to_slv(opcode_type, 16#08#),
      1901 => to_slv(opcode_type, 16#8C#),
      1902 => to_slv(opcode_type, 16#0B#),
      1903 => to_slv(opcode_type, 16#07#),
      1904 => to_slv(opcode_type, 16#07#),
      1905 => to_slv(opcode_type, 16#06#),
      1906 => to_slv(opcode_type, 16#10#),
      1907 => to_slv(opcode_type, 16#0F#),
      1908 => to_slv(opcode_type, 16#07#),
      1909 => to_slv(opcode_type, 16#0F#),
      1910 => to_slv(opcode_type, 16#0B#),
      1911 => to_slv(opcode_type, 16#07#),
      1912 => to_slv(opcode_type, 16#03#),
      1913 => to_slv(opcode_type, 16#76#),
      1914 => to_slv(opcode_type, 16#08#),
      1915 => to_slv(opcode_type, 16#0B#),
      1916 => to_slv(opcode_type, 16#0B#),
      1917 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#08#),
      1921 => to_slv(opcode_type, 16#06#),
      1922 => to_slv(opcode_type, 16#07#),
      1923 => to_slv(opcode_type, 16#09#),
      1924 => to_slv(opcode_type, 16#11#),
      1925 => to_slv(opcode_type, 16#0A#),
      1926 => to_slv(opcode_type, 16#02#),
      1927 => to_slv(opcode_type, 16#10#),
      1928 => to_slv(opcode_type, 16#07#),
      1929 => to_slv(opcode_type, 16#01#),
      1930 => to_slv(opcode_type, 16#0D#),
      1931 => to_slv(opcode_type, 16#06#),
      1932 => to_slv(opcode_type, 16#0A#),
      1933 => to_slv(opcode_type, 16#0C#),
      1934 => to_slv(opcode_type, 16#06#),
      1935 => to_slv(opcode_type, 16#09#),
      1936 => to_slv(opcode_type, 16#07#),
      1937 => to_slv(opcode_type, 16#0E#),
      1938 => to_slv(opcode_type, 16#0E#),
      1939 => to_slv(opcode_type, 16#09#),
      1940 => to_slv(opcode_type, 16#0F#),
      1941 => to_slv(opcode_type, 16#2E#),
      1942 => to_slv(opcode_type, 16#09#),
      1943 => to_slv(opcode_type, 16#09#),
      1944 => to_slv(opcode_type, 16#0C#),
      1945 => to_slv(opcode_type, 16#11#),
      1946 => to_slv(opcode_type, 16#06#),
      1947 => to_slv(opcode_type, 16#0C#),
      1948 => to_slv(opcode_type, 16#0E#),
      1949 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#07#),
      1953 => to_slv(opcode_type, 16#08#),
      1954 => to_slv(opcode_type, 16#06#),
      1955 => to_slv(opcode_type, 16#02#),
      1956 => to_slv(opcode_type, 16#10#),
      1957 => to_slv(opcode_type, 16#08#),
      1958 => to_slv(opcode_type, 16#0D#),
      1959 => to_slv(opcode_type, 16#0D#),
      1960 => to_slv(opcode_type, 16#08#),
      1961 => to_slv(opcode_type, 16#01#),
      1962 => to_slv(opcode_type, 16#0F#),
      1963 => to_slv(opcode_type, 16#08#),
      1964 => to_slv(opcode_type, 16#0D#),
      1965 => to_slv(opcode_type, 16#0E#),
      1966 => to_slv(opcode_type, 16#07#),
      1967 => to_slv(opcode_type, 16#09#),
      1968 => to_slv(opcode_type, 16#08#),
      1969 => to_slv(opcode_type, 16#11#),
      1970 => to_slv(opcode_type, 16#49#),
      1971 => to_slv(opcode_type, 16#06#),
      1972 => to_slv(opcode_type, 16#0A#),
      1973 => to_slv(opcode_type, 16#0E#),
      1974 => to_slv(opcode_type, 16#08#),
      1975 => to_slv(opcode_type, 16#08#),
      1976 => to_slv(opcode_type, 16#0C#),
      1977 => to_slv(opcode_type, 16#0F#),
      1978 => to_slv(opcode_type, 16#08#),
      1979 => to_slv(opcode_type, 16#0C#),
      1980 => to_slv(opcode_type, 16#0B#),
      1981 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#09#),
      1985 => to_slv(opcode_type, 16#07#),
      1986 => to_slv(opcode_type, 16#08#),
      1987 => to_slv(opcode_type, 16#08#),
      1988 => to_slv(opcode_type, 16#10#),
      1989 => to_slv(opcode_type, 16#11#),
      1990 => to_slv(opcode_type, 16#06#),
      1991 => to_slv(opcode_type, 16#0A#),
      1992 => to_slv(opcode_type, 16#0C#),
      1993 => to_slv(opcode_type, 16#07#),
      1994 => to_slv(opcode_type, 16#04#),
      1995 => to_slv(opcode_type, 16#0D#),
      1996 => to_slv(opcode_type, 16#04#),
      1997 => to_slv(opcode_type, 16#11#),
      1998 => to_slv(opcode_type, 16#08#),
      1999 => to_slv(opcode_type, 16#07#),
      2000 => to_slv(opcode_type, 16#06#),
      2001 => to_slv(opcode_type, 16#0A#),
      2002 => to_slv(opcode_type, 16#0E#),
      2003 => to_slv(opcode_type, 16#06#),
      2004 => to_slv(opcode_type, 16#0A#),
      2005 => to_slv(opcode_type, 16#0D#),
      2006 => to_slv(opcode_type, 16#09#),
      2007 => to_slv(opcode_type, 16#09#),
      2008 => to_slv(opcode_type, 16#0F#),
      2009 => to_slv(opcode_type, 16#10#),
      2010 => to_slv(opcode_type, 16#07#),
      2011 => to_slv(opcode_type, 16#0D#),
      2012 => to_slv(opcode_type, 16#0B#),
      2013 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#09#),
      2017 => to_slv(opcode_type, 16#08#),
      2018 => to_slv(opcode_type, 16#09#),
      2019 => to_slv(opcode_type, 16#01#),
      2020 => to_slv(opcode_type, 16#11#),
      2021 => to_slv(opcode_type, 16#09#),
      2022 => to_slv(opcode_type, 16#11#),
      2023 => to_slv(opcode_type, 16#0D#),
      2024 => to_slv(opcode_type, 16#07#),
      2025 => to_slv(opcode_type, 16#02#),
      2026 => to_slv(opcode_type, 16#0D#),
      2027 => to_slv(opcode_type, 16#08#),
      2028 => to_slv(opcode_type, 16#0F#),
      2029 => to_slv(opcode_type, 16#1E#),
      2030 => to_slv(opcode_type, 16#07#),
      2031 => to_slv(opcode_type, 16#09#),
      2032 => to_slv(opcode_type, 16#09#),
      2033 => to_slv(opcode_type, 16#0A#),
      2034 => to_slv(opcode_type, 16#0F#),
      2035 => to_slv(opcode_type, 16#06#),
      2036 => to_slv(opcode_type, 16#0E#),
      2037 => to_slv(opcode_type, 16#12#),
      2038 => to_slv(opcode_type, 16#07#),
      2039 => to_slv(opcode_type, 16#09#),
      2040 => to_slv(opcode_type, 16#0D#),
      2041 => to_slv(opcode_type, 16#0A#),
      2042 => to_slv(opcode_type, 16#06#),
      2043 => to_slv(opcode_type, 16#11#),
      2044 => to_slv(opcode_type, 16#0C#),
      2045 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#06#),
      2049 => to_slv(opcode_type, 16#07#),
      2050 => to_slv(opcode_type, 16#09#),
      2051 => to_slv(opcode_type, 16#03#),
      2052 => to_slv(opcode_type, 16#11#),
      2053 => to_slv(opcode_type, 16#02#),
      2054 => to_slv(opcode_type, 16#0F#),
      2055 => to_slv(opcode_type, 16#08#),
      2056 => to_slv(opcode_type, 16#06#),
      2057 => to_slv(opcode_type, 16#0A#),
      2058 => to_slv(opcode_type, 16#0E#),
      2059 => to_slv(opcode_type, 16#06#),
      2060 => to_slv(opcode_type, 16#0A#),
      2061 => to_slv(opcode_type, 16#11#),
      2062 => to_slv(opcode_type, 16#07#),
      2063 => to_slv(opcode_type, 16#07#),
      2064 => to_slv(opcode_type, 16#06#),
      2065 => to_slv(opcode_type, 16#0B#),
      2066 => to_slv(opcode_type, 16#0F#),
      2067 => to_slv(opcode_type, 16#09#),
      2068 => to_slv(opcode_type, 16#0A#),
      2069 => to_slv(opcode_type, 16#11#),
      2070 => to_slv(opcode_type, 16#07#),
      2071 => to_slv(opcode_type, 16#07#),
      2072 => to_slv(opcode_type, 16#0E#),
      2073 => to_slv(opcode_type, 16#0D#),
      2074 => to_slv(opcode_type, 16#06#),
      2075 => to_slv(opcode_type, 16#0D#),
      2076 => to_slv(opcode_type, 16#0D#),
      2077 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#09#),
      2081 => to_slv(opcode_type, 16#08#),
      2082 => to_slv(opcode_type, 16#08#),
      2083 => to_slv(opcode_type, 16#06#),
      2084 => to_slv(opcode_type, 16#0F#),
      2085 => to_slv(opcode_type, 16#0F#),
      2086 => to_slv(opcode_type, 16#05#),
      2087 => to_slv(opcode_type, 16#0D#),
      2088 => to_slv(opcode_type, 16#09#),
      2089 => to_slv(opcode_type, 16#02#),
      2090 => to_slv(opcode_type, 16#10#),
      2091 => to_slv(opcode_type, 16#07#),
      2092 => to_slv(opcode_type, 16#10#),
      2093 => to_slv(opcode_type, 16#0D#),
      2094 => to_slv(opcode_type, 16#09#),
      2095 => to_slv(opcode_type, 16#07#),
      2096 => to_slv(opcode_type, 16#09#),
      2097 => to_slv(opcode_type, 16#0C#),
      2098 => to_slv(opcode_type, 16#0C#),
      2099 => to_slv(opcode_type, 16#08#),
      2100 => to_slv(opcode_type, 16#53#),
      2101 => to_slv(opcode_type, 16#0B#),
      2102 => to_slv(opcode_type, 16#08#),
      2103 => to_slv(opcode_type, 16#06#),
      2104 => to_slv(opcode_type, 16#AD#),
      2105 => to_slv(opcode_type, 16#0D#),
      2106 => to_slv(opcode_type, 16#06#),
      2107 => to_slv(opcode_type, 16#10#),
      2108 => to_slv(opcode_type, 16#0F#),
      2109 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#06#),
      2113 => to_slv(opcode_type, 16#07#),
      2114 => to_slv(opcode_type, 16#06#),
      2115 => to_slv(opcode_type, 16#09#),
      2116 => to_slv(opcode_type, 16#11#),
      2117 => to_slv(opcode_type, 16#0A#),
      2118 => to_slv(opcode_type, 16#03#),
      2119 => to_slv(opcode_type, 16#0C#),
      2120 => to_slv(opcode_type, 16#06#),
      2121 => to_slv(opcode_type, 16#08#),
      2122 => to_slv(opcode_type, 16#10#),
      2123 => to_slv(opcode_type, 16#11#),
      2124 => to_slv(opcode_type, 16#03#),
      2125 => to_slv(opcode_type, 16#11#),
      2126 => to_slv(opcode_type, 16#08#),
      2127 => to_slv(opcode_type, 16#07#),
      2128 => to_slv(opcode_type, 16#06#),
      2129 => to_slv(opcode_type, 16#0F#),
      2130 => to_slv(opcode_type, 16#0A#),
      2131 => to_slv(opcode_type, 16#09#),
      2132 => to_slv(opcode_type, 16#0E#),
      2133 => to_slv(opcode_type, 16#0A#),
      2134 => to_slv(opcode_type, 16#09#),
      2135 => to_slv(opcode_type, 16#08#),
      2136 => to_slv(opcode_type, 16#0A#),
      2137 => to_slv(opcode_type, 16#0E#),
      2138 => to_slv(opcode_type, 16#09#),
      2139 => to_slv(opcode_type, 16#0D#),
      2140 => to_slv(opcode_type, 16#0B#),
      2141 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#09#),
      2146 => to_slv(opcode_type, 16#09#),
      2147 => to_slv(opcode_type, 16#08#),
      2148 => to_slv(opcode_type, 16#9B#),
      2149 => to_slv(opcode_type, 16#E4#),
      2150 => to_slv(opcode_type, 16#07#),
      2151 => to_slv(opcode_type, 16#0E#),
      2152 => to_slv(opcode_type, 16#0D#),
      2153 => to_slv(opcode_type, 16#08#),
      2154 => to_slv(opcode_type, 16#07#),
      2155 => to_slv(opcode_type, 16#10#),
      2156 => to_slv(opcode_type, 16#0F#),
      2157 => to_slv(opcode_type, 16#01#),
      2158 => to_slv(opcode_type, 16#0C#),
      2159 => to_slv(opcode_type, 16#07#),
      2160 => to_slv(opcode_type, 16#06#),
      2161 => to_slv(opcode_type, 16#07#),
      2162 => to_slv(opcode_type, 16#0C#),
      2163 => to_slv(opcode_type, 16#0D#),
      2164 => to_slv(opcode_type, 16#01#),
      2165 => to_slv(opcode_type, 16#4A#),
      2166 => to_slv(opcode_type, 16#07#),
      2167 => to_slv(opcode_type, 16#08#),
      2168 => to_slv(opcode_type, 16#0A#),
      2169 => to_slv(opcode_type, 16#0D#),
      2170 => to_slv(opcode_type, 16#08#),
      2171 => to_slv(opcode_type, 16#0F#),
      2172 => to_slv(opcode_type, 16#6C#),
      2173 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#08#),
      2177 => to_slv(opcode_type, 16#09#),
      2178 => to_slv(opcode_type, 16#06#),
      2179 => to_slv(opcode_type, 16#02#),
      2180 => to_slv(opcode_type, 16#0C#),
      2181 => to_slv(opcode_type, 16#05#),
      2182 => to_slv(opcode_type, 16#0A#),
      2183 => to_slv(opcode_type, 16#07#),
      2184 => to_slv(opcode_type, 16#06#),
      2185 => to_slv(opcode_type, 16#0C#),
      2186 => to_slv(opcode_type, 16#11#),
      2187 => to_slv(opcode_type, 16#08#),
      2188 => to_slv(opcode_type, 16#0B#),
      2189 => to_slv(opcode_type, 16#0C#),
      2190 => to_slv(opcode_type, 16#09#),
      2191 => to_slv(opcode_type, 16#09#),
      2192 => to_slv(opcode_type, 16#08#),
      2193 => to_slv(opcode_type, 16#0E#),
      2194 => to_slv(opcode_type, 16#F4#),
      2195 => to_slv(opcode_type, 16#07#),
      2196 => to_slv(opcode_type, 16#A6#),
      2197 => to_slv(opcode_type, 16#0F#),
      2198 => to_slv(opcode_type, 16#08#),
      2199 => to_slv(opcode_type, 16#08#),
      2200 => to_slv(opcode_type, 16#0D#),
      2201 => to_slv(opcode_type, 16#0C#),
      2202 => to_slv(opcode_type, 16#06#),
      2203 => to_slv(opcode_type, 16#11#),
      2204 => to_slv(opcode_type, 16#0F#),
      2205 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#08#),
      2209 => to_slv(opcode_type, 16#08#),
      2210 => to_slv(opcode_type, 16#09#),
      2211 => to_slv(opcode_type, 16#04#),
      2212 => to_slv(opcode_type, 16#0C#),
      2213 => to_slv(opcode_type, 16#03#),
      2214 => to_slv(opcode_type, 16#0A#),
      2215 => to_slv(opcode_type, 16#06#),
      2216 => to_slv(opcode_type, 16#07#),
      2217 => to_slv(opcode_type, 16#0E#),
      2218 => to_slv(opcode_type, 16#0A#),
      2219 => to_slv(opcode_type, 16#06#),
      2220 => to_slv(opcode_type, 16#0A#),
      2221 => to_slv(opcode_type, 16#0E#),
      2222 => to_slv(opcode_type, 16#09#),
      2223 => to_slv(opcode_type, 16#08#),
      2224 => to_slv(opcode_type, 16#06#),
      2225 => to_slv(opcode_type, 16#11#),
      2226 => to_slv(opcode_type, 16#0A#),
      2227 => to_slv(opcode_type, 16#08#),
      2228 => to_slv(opcode_type, 16#11#),
      2229 => to_slv(opcode_type, 16#0C#),
      2230 => to_slv(opcode_type, 16#09#),
      2231 => to_slv(opcode_type, 16#08#),
      2232 => to_slv(opcode_type, 16#0B#),
      2233 => to_slv(opcode_type, 16#0E#),
      2234 => to_slv(opcode_type, 16#06#),
      2235 => to_slv(opcode_type, 16#0E#),
      2236 => to_slv(opcode_type, 16#CC#),
      2237 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#09#),
      2242 => to_slv(opcode_type, 16#07#),
      2243 => to_slv(opcode_type, 16#03#),
      2244 => to_slv(opcode_type, 16#0E#),
      2245 => to_slv(opcode_type, 16#04#),
      2246 => to_slv(opcode_type, 16#0A#),
      2247 => to_slv(opcode_type, 16#08#),
      2248 => to_slv(opcode_type, 16#07#),
      2249 => to_slv(opcode_type, 16#11#),
      2250 => to_slv(opcode_type, 16#0A#),
      2251 => to_slv(opcode_type, 16#08#),
      2252 => to_slv(opcode_type, 16#0A#),
      2253 => to_slv(opcode_type, 16#0D#),
      2254 => to_slv(opcode_type, 16#07#),
      2255 => to_slv(opcode_type, 16#08#),
      2256 => to_slv(opcode_type, 16#08#),
      2257 => to_slv(opcode_type, 16#0E#),
      2258 => to_slv(opcode_type, 16#11#),
      2259 => to_slv(opcode_type, 16#09#),
      2260 => to_slv(opcode_type, 16#10#),
      2261 => to_slv(opcode_type, 16#0A#),
      2262 => to_slv(opcode_type, 16#08#),
      2263 => to_slv(opcode_type, 16#09#),
      2264 => to_slv(opcode_type, 16#0F#),
      2265 => to_slv(opcode_type, 16#2C#),
      2266 => to_slv(opcode_type, 16#09#),
      2267 => to_slv(opcode_type, 16#11#),
      2268 => to_slv(opcode_type, 16#0E#),
      2269 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#06#),
      2273 => to_slv(opcode_type, 16#07#),
      2274 => to_slv(opcode_type, 16#08#),
      2275 => to_slv(opcode_type, 16#09#),
      2276 => to_slv(opcode_type, 16#5A#),
      2277 => to_slv(opcode_type, 16#0D#),
      2278 => to_slv(opcode_type, 16#04#),
      2279 => to_slv(opcode_type, 16#10#),
      2280 => to_slv(opcode_type, 16#06#),
      2281 => to_slv(opcode_type, 16#04#),
      2282 => to_slv(opcode_type, 16#0F#),
      2283 => to_slv(opcode_type, 16#07#),
      2284 => to_slv(opcode_type, 16#0B#),
      2285 => to_slv(opcode_type, 16#11#),
      2286 => to_slv(opcode_type, 16#08#),
      2287 => to_slv(opcode_type, 16#06#),
      2288 => to_slv(opcode_type, 16#09#),
      2289 => to_slv(opcode_type, 16#CE#),
      2290 => to_slv(opcode_type, 16#10#),
      2291 => to_slv(opcode_type, 16#09#),
      2292 => to_slv(opcode_type, 16#0C#),
      2293 => to_slv(opcode_type, 16#32#),
      2294 => to_slv(opcode_type, 16#08#),
      2295 => to_slv(opcode_type, 16#07#),
      2296 => to_slv(opcode_type, 16#0C#),
      2297 => to_slv(opcode_type, 16#10#),
      2298 => to_slv(opcode_type, 16#09#),
      2299 => to_slv(opcode_type, 16#0D#),
      2300 => to_slv(opcode_type, 16#0D#),
      2301 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#07#),
      2305 => to_slv(opcode_type, 16#07#),
      2306 => to_slv(opcode_type, 16#06#),
      2307 => to_slv(opcode_type, 16#07#),
      2308 => to_slv(opcode_type, 16#0A#),
      2309 => to_slv(opcode_type, 16#0A#),
      2310 => to_slv(opcode_type, 16#05#),
      2311 => to_slv(opcode_type, 16#0F#),
      2312 => to_slv(opcode_type, 16#08#),
      2313 => to_slv(opcode_type, 16#08#),
      2314 => to_slv(opcode_type, 16#0D#),
      2315 => to_slv(opcode_type, 16#10#),
      2316 => to_slv(opcode_type, 16#02#),
      2317 => to_slv(opcode_type, 16#0F#),
      2318 => to_slv(opcode_type, 16#08#),
      2319 => to_slv(opcode_type, 16#06#),
      2320 => to_slv(opcode_type, 16#06#),
      2321 => to_slv(opcode_type, 16#0B#),
      2322 => to_slv(opcode_type, 16#10#),
      2323 => to_slv(opcode_type, 16#09#),
      2324 => to_slv(opcode_type, 16#0B#),
      2325 => to_slv(opcode_type, 16#0C#),
      2326 => to_slv(opcode_type, 16#09#),
      2327 => to_slv(opcode_type, 16#06#),
      2328 => to_slv(opcode_type, 16#11#),
      2329 => to_slv(opcode_type, 16#0C#),
      2330 => to_slv(opcode_type, 16#07#),
      2331 => to_slv(opcode_type, 16#9F#),
      2332 => to_slv(opcode_type, 16#0A#),
      2333 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#06#),
      2337 => to_slv(opcode_type, 16#08#),
      2338 => to_slv(opcode_type, 16#06#),
      2339 => to_slv(opcode_type, 16#06#),
      2340 => to_slv(opcode_type, 16#0B#),
      2341 => to_slv(opcode_type, 16#0F#),
      2342 => to_slv(opcode_type, 16#07#),
      2343 => to_slv(opcode_type, 16#0E#),
      2344 => to_slv(opcode_type, 16#0B#),
      2345 => to_slv(opcode_type, 16#08#),
      2346 => to_slv(opcode_type, 16#04#),
      2347 => to_slv(opcode_type, 16#67#),
      2348 => to_slv(opcode_type, 16#01#),
      2349 => to_slv(opcode_type, 16#0B#),
      2350 => to_slv(opcode_type, 16#08#),
      2351 => to_slv(opcode_type, 16#06#),
      2352 => to_slv(opcode_type, 16#09#),
      2353 => to_slv(opcode_type, 16#0B#),
      2354 => to_slv(opcode_type, 16#0C#),
      2355 => to_slv(opcode_type, 16#06#),
      2356 => to_slv(opcode_type, 16#0D#),
      2357 => to_slv(opcode_type, 16#0D#),
      2358 => to_slv(opcode_type, 16#09#),
      2359 => to_slv(opcode_type, 16#09#),
      2360 => to_slv(opcode_type, 16#11#),
      2361 => to_slv(opcode_type, 16#0F#),
      2362 => to_slv(opcode_type, 16#07#),
      2363 => to_slv(opcode_type, 16#11#),
      2364 => to_slv(opcode_type, 16#0F#),
      2365 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#07#),
      2369 => to_slv(opcode_type, 16#08#),
      2370 => to_slv(opcode_type, 16#08#),
      2371 => to_slv(opcode_type, 16#05#),
      2372 => to_slv(opcode_type, 16#0C#),
      2373 => to_slv(opcode_type, 16#05#),
      2374 => to_slv(opcode_type, 16#3A#),
      2375 => to_slv(opcode_type, 16#08#),
      2376 => to_slv(opcode_type, 16#08#),
      2377 => to_slv(opcode_type, 16#0F#),
      2378 => to_slv(opcode_type, 16#0C#),
      2379 => to_slv(opcode_type, 16#09#),
      2380 => to_slv(opcode_type, 16#10#),
      2381 => to_slv(opcode_type, 16#0D#),
      2382 => to_slv(opcode_type, 16#06#),
      2383 => to_slv(opcode_type, 16#09#),
      2384 => to_slv(opcode_type, 16#07#),
      2385 => to_slv(opcode_type, 16#F5#),
      2386 => to_slv(opcode_type, 16#11#),
      2387 => to_slv(opcode_type, 16#07#),
      2388 => to_slv(opcode_type, 16#0C#),
      2389 => to_slv(opcode_type, 16#0B#),
      2390 => to_slv(opcode_type, 16#06#),
      2391 => to_slv(opcode_type, 16#09#),
      2392 => to_slv(opcode_type, 16#0E#),
      2393 => to_slv(opcode_type, 16#0F#),
      2394 => to_slv(opcode_type, 16#06#),
      2395 => to_slv(opcode_type, 16#0B#),
      2396 => to_slv(opcode_type, 16#0D#),
      2397 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#07#),
      2401 => to_slv(opcode_type, 16#08#),
      2402 => to_slv(opcode_type, 16#08#),
      2403 => to_slv(opcode_type, 16#05#),
      2404 => to_slv(opcode_type, 16#0B#),
      2405 => to_slv(opcode_type, 16#05#),
      2406 => to_slv(opcode_type, 16#0C#),
      2407 => to_slv(opcode_type, 16#07#),
      2408 => to_slv(opcode_type, 16#07#),
      2409 => to_slv(opcode_type, 16#0D#),
      2410 => to_slv(opcode_type, 16#10#),
      2411 => to_slv(opcode_type, 16#08#),
      2412 => to_slv(opcode_type, 16#0A#),
      2413 => to_slv(opcode_type, 16#0E#),
      2414 => to_slv(opcode_type, 16#09#),
      2415 => to_slv(opcode_type, 16#09#),
      2416 => to_slv(opcode_type, 16#08#),
      2417 => to_slv(opcode_type, 16#0F#),
      2418 => to_slv(opcode_type, 16#0A#),
      2419 => to_slv(opcode_type, 16#07#),
      2420 => to_slv(opcode_type, 16#10#),
      2421 => to_slv(opcode_type, 16#6D#),
      2422 => to_slv(opcode_type, 16#06#),
      2423 => to_slv(opcode_type, 16#08#),
      2424 => to_slv(opcode_type, 16#0B#),
      2425 => to_slv(opcode_type, 16#0D#),
      2426 => to_slv(opcode_type, 16#08#),
      2427 => to_slv(opcode_type, 16#0E#),
      2428 => to_slv(opcode_type, 16#0D#),
      2429 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#07#),
      2433 => to_slv(opcode_type, 16#08#),
      2434 => to_slv(opcode_type, 16#07#),
      2435 => to_slv(opcode_type, 16#04#),
      2436 => to_slv(opcode_type, 16#0F#),
      2437 => to_slv(opcode_type, 16#04#),
      2438 => to_slv(opcode_type, 16#0F#),
      2439 => to_slv(opcode_type, 16#07#),
      2440 => to_slv(opcode_type, 16#08#),
      2441 => to_slv(opcode_type, 16#0D#),
      2442 => to_slv(opcode_type, 16#0B#),
      2443 => to_slv(opcode_type, 16#08#),
      2444 => to_slv(opcode_type, 16#0E#),
      2445 => to_slv(opcode_type, 16#0E#),
      2446 => to_slv(opcode_type, 16#08#),
      2447 => to_slv(opcode_type, 16#09#),
      2448 => to_slv(opcode_type, 16#07#),
      2449 => to_slv(opcode_type, 16#0B#),
      2450 => to_slv(opcode_type, 16#11#),
      2451 => to_slv(opcode_type, 16#06#),
      2452 => to_slv(opcode_type, 16#10#),
      2453 => to_slv(opcode_type, 16#0C#),
      2454 => to_slv(opcode_type, 16#08#),
      2455 => to_slv(opcode_type, 16#08#),
      2456 => to_slv(opcode_type, 16#0C#),
      2457 => to_slv(opcode_type, 16#0E#),
      2458 => to_slv(opcode_type, 16#09#),
      2459 => to_slv(opcode_type, 16#10#),
      2460 => to_slv(opcode_type, 16#FE#),
      2461 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#09#),
      2465 => to_slv(opcode_type, 16#09#),
      2466 => to_slv(opcode_type, 16#08#),
      2467 => to_slv(opcode_type, 16#03#),
      2468 => to_slv(opcode_type, 16#10#),
      2469 => to_slv(opcode_type, 16#05#),
      2470 => to_slv(opcode_type, 16#0B#),
      2471 => to_slv(opcode_type, 16#08#),
      2472 => to_slv(opcode_type, 16#08#),
      2473 => to_slv(opcode_type, 16#11#),
      2474 => to_slv(opcode_type, 16#D0#),
      2475 => to_slv(opcode_type, 16#09#),
      2476 => to_slv(opcode_type, 16#0D#),
      2477 => to_slv(opcode_type, 16#0A#),
      2478 => to_slv(opcode_type, 16#09#),
      2479 => to_slv(opcode_type, 16#09#),
      2480 => to_slv(opcode_type, 16#09#),
      2481 => to_slv(opcode_type, 16#0F#),
      2482 => to_slv(opcode_type, 16#0E#),
      2483 => to_slv(opcode_type, 16#06#),
      2484 => to_slv(opcode_type, 16#10#),
      2485 => to_slv(opcode_type, 16#11#),
      2486 => to_slv(opcode_type, 16#07#),
      2487 => to_slv(opcode_type, 16#07#),
      2488 => to_slv(opcode_type, 16#0F#),
      2489 => to_slv(opcode_type, 16#0F#),
      2490 => to_slv(opcode_type, 16#06#),
      2491 => to_slv(opcode_type, 16#40#),
      2492 => to_slv(opcode_type, 16#0E#),
      2493 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#06#),
      2497 => to_slv(opcode_type, 16#06#),
      2498 => to_slv(opcode_type, 16#09#),
      2499 => to_slv(opcode_type, 16#09#),
      2500 => to_slv(opcode_type, 16#0F#),
      2501 => to_slv(opcode_type, 16#0D#),
      2502 => to_slv(opcode_type, 16#05#),
      2503 => to_slv(opcode_type, 16#A3#),
      2504 => to_slv(opcode_type, 16#09#),
      2505 => to_slv(opcode_type, 16#07#),
      2506 => to_slv(opcode_type, 16#0D#),
      2507 => to_slv(opcode_type, 16#0B#),
      2508 => to_slv(opcode_type, 16#06#),
      2509 => to_slv(opcode_type, 16#0A#),
      2510 => to_slv(opcode_type, 16#0B#),
      2511 => to_slv(opcode_type, 16#07#),
      2512 => to_slv(opcode_type, 16#08#),
      2513 => to_slv(opcode_type, 16#06#),
      2514 => to_slv(opcode_type, 16#0B#),
      2515 => to_slv(opcode_type, 16#0A#),
      2516 => to_slv(opcode_type, 16#03#),
      2517 => to_slv(opcode_type, 16#0A#),
      2518 => to_slv(opcode_type, 16#07#),
      2519 => to_slv(opcode_type, 16#07#),
      2520 => to_slv(opcode_type, 16#0C#),
      2521 => to_slv(opcode_type, 16#0F#),
      2522 => to_slv(opcode_type, 16#07#),
      2523 => to_slv(opcode_type, 16#0F#),
      2524 => to_slv(opcode_type, 16#0C#),
      2525 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#07#),
      2529 => to_slv(opcode_type, 16#08#),
      2530 => to_slv(opcode_type, 16#06#),
      2531 => to_slv(opcode_type, 16#09#),
      2532 => to_slv(opcode_type, 16#10#),
      2533 => to_slv(opcode_type, 16#0F#),
      2534 => to_slv(opcode_type, 16#04#),
      2535 => to_slv(opcode_type, 16#0E#),
      2536 => to_slv(opcode_type, 16#07#),
      2537 => to_slv(opcode_type, 16#06#),
      2538 => to_slv(opcode_type, 16#10#),
      2539 => to_slv(opcode_type, 16#11#),
      2540 => to_slv(opcode_type, 16#04#),
      2541 => to_slv(opcode_type, 16#11#),
      2542 => to_slv(opcode_type, 16#07#),
      2543 => to_slv(opcode_type, 16#06#),
      2544 => to_slv(opcode_type, 16#07#),
      2545 => to_slv(opcode_type, 16#B0#),
      2546 => to_slv(opcode_type, 16#0A#),
      2547 => to_slv(opcode_type, 16#07#),
      2548 => to_slv(opcode_type, 16#0F#),
      2549 => to_slv(opcode_type, 16#0F#),
      2550 => to_slv(opcode_type, 16#08#),
      2551 => to_slv(opcode_type, 16#08#),
      2552 => to_slv(opcode_type, 16#0A#),
      2553 => to_slv(opcode_type, 16#11#),
      2554 => to_slv(opcode_type, 16#07#),
      2555 => to_slv(opcode_type, 16#11#),
      2556 => to_slv(opcode_type, 16#95#),
      2557 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#07#),
      2561 => to_slv(opcode_type, 16#09#),
      2562 => to_slv(opcode_type, 16#08#),
      2563 => to_slv(opcode_type, 16#07#),
      2564 => to_slv(opcode_type, 16#0D#),
      2565 => to_slv(opcode_type, 16#0B#),
      2566 => to_slv(opcode_type, 16#07#),
      2567 => to_slv(opcode_type, 16#0F#),
      2568 => to_slv(opcode_type, 16#11#),
      2569 => to_slv(opcode_type, 16#06#),
      2570 => to_slv(opcode_type, 16#04#),
      2571 => to_slv(opcode_type, 16#FF#),
      2572 => to_slv(opcode_type, 16#03#),
      2573 => to_slv(opcode_type, 16#9E#),
      2574 => to_slv(opcode_type, 16#07#),
      2575 => to_slv(opcode_type, 16#08#),
      2576 => to_slv(opcode_type, 16#06#),
      2577 => to_slv(opcode_type, 16#10#),
      2578 => to_slv(opcode_type, 16#0D#),
      2579 => to_slv(opcode_type, 16#07#),
      2580 => to_slv(opcode_type, 16#0A#),
      2581 => to_slv(opcode_type, 16#0A#),
      2582 => to_slv(opcode_type, 16#07#),
      2583 => to_slv(opcode_type, 16#09#),
      2584 => to_slv(opcode_type, 16#54#),
      2585 => to_slv(opcode_type, 16#0F#),
      2586 => to_slv(opcode_type, 16#08#),
      2587 => to_slv(opcode_type, 16#11#),
      2588 => to_slv(opcode_type, 16#0C#),
      2589 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#09#),
      2593 => to_slv(opcode_type, 16#07#),
      2594 => to_slv(opcode_type, 16#09#),
      2595 => to_slv(opcode_type, 16#09#),
      2596 => to_slv(opcode_type, 16#10#),
      2597 => to_slv(opcode_type, 16#0A#),
      2598 => to_slv(opcode_type, 16#02#),
      2599 => to_slv(opcode_type, 16#0F#),
      2600 => to_slv(opcode_type, 16#08#),
      2601 => to_slv(opcode_type, 16#09#),
      2602 => to_slv(opcode_type, 16#0D#),
      2603 => to_slv(opcode_type, 16#0A#),
      2604 => to_slv(opcode_type, 16#06#),
      2605 => to_slv(opcode_type, 16#EC#),
      2606 => to_slv(opcode_type, 16#0A#),
      2607 => to_slv(opcode_type, 16#07#),
      2608 => to_slv(opcode_type, 16#09#),
      2609 => to_slv(opcode_type, 16#05#),
      2610 => to_slv(opcode_type, 16#0C#),
      2611 => to_slv(opcode_type, 16#06#),
      2612 => to_slv(opcode_type, 16#10#),
      2613 => to_slv(opcode_type, 16#0C#),
      2614 => to_slv(opcode_type, 16#09#),
      2615 => to_slv(opcode_type, 16#06#),
      2616 => to_slv(opcode_type, 16#0C#),
      2617 => to_slv(opcode_type, 16#0C#),
      2618 => to_slv(opcode_type, 16#06#),
      2619 => to_slv(opcode_type, 16#10#),
      2620 => to_slv(opcode_type, 16#0A#),
      2621 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#09#),
      2625 => to_slv(opcode_type, 16#06#),
      2626 => to_slv(opcode_type, 16#07#),
      2627 => to_slv(opcode_type, 16#03#),
      2628 => to_slv(opcode_type, 16#0F#),
      2629 => to_slv(opcode_type, 16#08#),
      2630 => to_slv(opcode_type, 16#68#),
      2631 => to_slv(opcode_type, 16#0D#),
      2632 => to_slv(opcode_type, 16#08#),
      2633 => to_slv(opcode_type, 16#01#),
      2634 => to_slv(opcode_type, 16#5F#),
      2635 => to_slv(opcode_type, 16#09#),
      2636 => to_slv(opcode_type, 16#0C#),
      2637 => to_slv(opcode_type, 16#0B#),
      2638 => to_slv(opcode_type, 16#07#),
      2639 => to_slv(opcode_type, 16#06#),
      2640 => to_slv(opcode_type, 16#06#),
      2641 => to_slv(opcode_type, 16#0D#),
      2642 => to_slv(opcode_type, 16#0E#),
      2643 => to_slv(opcode_type, 16#06#),
      2644 => to_slv(opcode_type, 16#10#),
      2645 => to_slv(opcode_type, 16#E4#),
      2646 => to_slv(opcode_type, 16#08#),
      2647 => to_slv(opcode_type, 16#07#),
      2648 => to_slv(opcode_type, 16#8C#),
      2649 => to_slv(opcode_type, 16#0A#),
      2650 => to_slv(opcode_type, 16#06#),
      2651 => to_slv(opcode_type, 16#11#),
      2652 => to_slv(opcode_type, 16#11#),
      2653 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#09#),
      2657 => to_slv(opcode_type, 16#07#),
      2658 => to_slv(opcode_type, 16#08#),
      2659 => to_slv(opcode_type, 16#05#),
      2660 => to_slv(opcode_type, 16#0A#),
      2661 => to_slv(opcode_type, 16#09#),
      2662 => to_slv(opcode_type, 16#0B#),
      2663 => to_slv(opcode_type, 16#11#),
      2664 => to_slv(opcode_type, 16#09#),
      2665 => to_slv(opcode_type, 16#06#),
      2666 => to_slv(opcode_type, 16#0C#),
      2667 => to_slv(opcode_type, 16#10#),
      2668 => to_slv(opcode_type, 16#09#),
      2669 => to_slv(opcode_type, 16#0F#),
      2670 => to_slv(opcode_type, 16#10#),
      2671 => to_slv(opcode_type, 16#07#),
      2672 => to_slv(opcode_type, 16#06#),
      2673 => to_slv(opcode_type, 16#04#),
      2674 => to_slv(opcode_type, 16#11#),
      2675 => to_slv(opcode_type, 16#09#),
      2676 => to_slv(opcode_type, 16#0E#),
      2677 => to_slv(opcode_type, 16#0C#),
      2678 => to_slv(opcode_type, 16#08#),
      2679 => to_slv(opcode_type, 16#09#),
      2680 => to_slv(opcode_type, 16#0F#),
      2681 => to_slv(opcode_type, 16#0B#),
      2682 => to_slv(opcode_type, 16#07#),
      2683 => to_slv(opcode_type, 16#0E#),
      2684 => to_slv(opcode_type, 16#0B#),
      2685 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#06#),
      2689 => to_slv(opcode_type, 16#07#),
      2690 => to_slv(opcode_type, 16#08#),
      2691 => to_slv(opcode_type, 16#05#),
      2692 => to_slv(opcode_type, 16#0C#),
      2693 => to_slv(opcode_type, 16#02#),
      2694 => to_slv(opcode_type, 16#0F#),
      2695 => to_slv(opcode_type, 16#06#),
      2696 => to_slv(opcode_type, 16#09#),
      2697 => to_slv(opcode_type, 16#0C#),
      2698 => to_slv(opcode_type, 16#0E#),
      2699 => to_slv(opcode_type, 16#06#),
      2700 => to_slv(opcode_type, 16#10#),
      2701 => to_slv(opcode_type, 16#0F#),
      2702 => to_slv(opcode_type, 16#08#),
      2703 => to_slv(opcode_type, 16#06#),
      2704 => to_slv(opcode_type, 16#06#),
      2705 => to_slv(opcode_type, 16#FE#),
      2706 => to_slv(opcode_type, 16#0D#),
      2707 => to_slv(opcode_type, 16#08#),
      2708 => to_slv(opcode_type, 16#0C#),
      2709 => to_slv(opcode_type, 16#0F#),
      2710 => to_slv(opcode_type, 16#06#),
      2711 => to_slv(opcode_type, 16#06#),
      2712 => to_slv(opcode_type, 16#0A#),
      2713 => to_slv(opcode_type, 16#0D#),
      2714 => to_slv(opcode_type, 16#06#),
      2715 => to_slv(opcode_type, 16#0A#),
      2716 => to_slv(opcode_type, 16#0C#),
      2717 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#06#),
      2721 => to_slv(opcode_type, 16#09#),
      2722 => to_slv(opcode_type, 16#06#),
      2723 => to_slv(opcode_type, 16#04#),
      2724 => to_slv(opcode_type, 16#0D#),
      2725 => to_slv(opcode_type, 16#01#),
      2726 => to_slv(opcode_type, 16#83#),
      2727 => to_slv(opcode_type, 16#07#),
      2728 => to_slv(opcode_type, 16#09#),
      2729 => to_slv(opcode_type, 16#0C#),
      2730 => to_slv(opcode_type, 16#0C#),
      2731 => to_slv(opcode_type, 16#09#),
      2732 => to_slv(opcode_type, 16#11#),
      2733 => to_slv(opcode_type, 16#0B#),
      2734 => to_slv(opcode_type, 16#08#),
      2735 => to_slv(opcode_type, 16#09#),
      2736 => to_slv(opcode_type, 16#07#),
      2737 => to_slv(opcode_type, 16#0E#),
      2738 => to_slv(opcode_type, 16#0E#),
      2739 => to_slv(opcode_type, 16#06#),
      2740 => to_slv(opcode_type, 16#0E#),
      2741 => to_slv(opcode_type, 16#0E#),
      2742 => to_slv(opcode_type, 16#07#),
      2743 => to_slv(opcode_type, 16#07#),
      2744 => to_slv(opcode_type, 16#0C#),
      2745 => to_slv(opcode_type, 16#0A#),
      2746 => to_slv(opcode_type, 16#07#),
      2747 => to_slv(opcode_type, 16#10#),
      2748 => to_slv(opcode_type, 16#11#),
      2749 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#06#),
      2753 => to_slv(opcode_type, 16#09#),
      2754 => to_slv(opcode_type, 16#08#),
      2755 => to_slv(opcode_type, 16#09#),
      2756 => to_slv(opcode_type, 16#0E#),
      2757 => to_slv(opcode_type, 16#0B#),
      2758 => to_slv(opcode_type, 16#06#),
      2759 => to_slv(opcode_type, 16#11#),
      2760 => to_slv(opcode_type, 16#11#),
      2761 => to_slv(opcode_type, 16#09#),
      2762 => to_slv(opcode_type, 16#08#),
      2763 => to_slv(opcode_type, 16#0A#),
      2764 => to_slv(opcode_type, 16#11#),
      2765 => to_slv(opcode_type, 16#03#),
      2766 => to_slv(opcode_type, 16#0A#),
      2767 => to_slv(opcode_type, 16#09#),
      2768 => to_slv(opcode_type, 16#09#),
      2769 => to_slv(opcode_type, 16#07#),
      2770 => to_slv(opcode_type, 16#0F#),
      2771 => to_slv(opcode_type, 16#CC#),
      2772 => to_slv(opcode_type, 16#06#),
      2773 => to_slv(opcode_type, 16#0B#),
      2774 => to_slv(opcode_type, 16#0C#),
      2775 => to_slv(opcode_type, 16#06#),
      2776 => to_slv(opcode_type, 16#01#),
      2777 => to_slv(opcode_type, 16#0F#),
      2778 => to_slv(opcode_type, 16#08#),
      2779 => to_slv(opcode_type, 16#11#),
      2780 => to_slv(opcode_type, 16#0E#),
      2781 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#09#),
      2785 => to_slv(opcode_type, 16#09#),
      2786 => to_slv(opcode_type, 16#08#),
      2787 => to_slv(opcode_type, 16#01#),
      2788 => to_slv(opcode_type, 16#11#),
      2789 => to_slv(opcode_type, 16#03#),
      2790 => to_slv(opcode_type, 16#0D#),
      2791 => to_slv(opcode_type, 16#08#),
      2792 => to_slv(opcode_type, 16#08#),
      2793 => to_slv(opcode_type, 16#0F#),
      2794 => to_slv(opcode_type, 16#11#),
      2795 => to_slv(opcode_type, 16#06#),
      2796 => to_slv(opcode_type, 16#11#),
      2797 => to_slv(opcode_type, 16#11#),
      2798 => to_slv(opcode_type, 16#07#),
      2799 => to_slv(opcode_type, 16#09#),
      2800 => to_slv(opcode_type, 16#08#),
      2801 => to_slv(opcode_type, 16#0B#),
      2802 => to_slv(opcode_type, 16#10#),
      2803 => to_slv(opcode_type, 16#07#),
      2804 => to_slv(opcode_type, 16#10#),
      2805 => to_slv(opcode_type, 16#11#),
      2806 => to_slv(opcode_type, 16#07#),
      2807 => to_slv(opcode_type, 16#06#),
      2808 => to_slv(opcode_type, 16#0C#),
      2809 => to_slv(opcode_type, 16#43#),
      2810 => to_slv(opcode_type, 16#07#),
      2811 => to_slv(opcode_type, 16#10#),
      2812 => to_slv(opcode_type, 16#11#),
      2813 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#09#),
      2817 => to_slv(opcode_type, 16#06#),
      2818 => to_slv(opcode_type, 16#08#),
      2819 => to_slv(opcode_type, 16#04#),
      2820 => to_slv(opcode_type, 16#0D#),
      2821 => to_slv(opcode_type, 16#08#),
      2822 => to_slv(opcode_type, 16#0C#),
      2823 => to_slv(opcode_type, 16#11#),
      2824 => to_slv(opcode_type, 16#08#),
      2825 => to_slv(opcode_type, 16#01#),
      2826 => to_slv(opcode_type, 16#0A#),
      2827 => to_slv(opcode_type, 16#08#),
      2828 => to_slv(opcode_type, 16#0F#),
      2829 => to_slv(opcode_type, 16#10#),
      2830 => to_slv(opcode_type, 16#06#),
      2831 => to_slv(opcode_type, 16#09#),
      2832 => to_slv(opcode_type, 16#09#),
      2833 => to_slv(opcode_type, 16#0C#),
      2834 => to_slv(opcode_type, 16#0D#),
      2835 => to_slv(opcode_type, 16#07#),
      2836 => to_slv(opcode_type, 16#0B#),
      2837 => to_slv(opcode_type, 16#F6#),
      2838 => to_slv(opcode_type, 16#08#),
      2839 => to_slv(opcode_type, 16#09#),
      2840 => to_slv(opcode_type, 16#3A#),
      2841 => to_slv(opcode_type, 16#0B#),
      2842 => to_slv(opcode_type, 16#09#),
      2843 => to_slv(opcode_type, 16#0C#),
      2844 => to_slv(opcode_type, 16#0C#),
      2845 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#06#),
      2849 => to_slv(opcode_type, 16#07#),
      2850 => to_slv(opcode_type, 16#06#),
      2851 => to_slv(opcode_type, 16#07#),
      2852 => to_slv(opcode_type, 16#0F#),
      2853 => to_slv(opcode_type, 16#0C#),
      2854 => to_slv(opcode_type, 16#03#),
      2855 => to_slv(opcode_type, 16#0E#),
      2856 => to_slv(opcode_type, 16#09#),
      2857 => to_slv(opcode_type, 16#09#),
      2858 => to_slv(opcode_type, 16#0E#),
      2859 => to_slv(opcode_type, 16#0D#),
      2860 => to_slv(opcode_type, 16#06#),
      2861 => to_slv(opcode_type, 16#0E#),
      2862 => to_slv(opcode_type, 16#10#),
      2863 => to_slv(opcode_type, 16#06#),
      2864 => to_slv(opcode_type, 16#06#),
      2865 => to_slv(opcode_type, 16#01#),
      2866 => to_slv(opcode_type, 16#0B#),
      2867 => to_slv(opcode_type, 16#07#),
      2868 => to_slv(opcode_type, 16#0D#),
      2869 => to_slv(opcode_type, 16#0E#),
      2870 => to_slv(opcode_type, 16#06#),
      2871 => to_slv(opcode_type, 16#09#),
      2872 => to_slv(opcode_type, 16#0C#),
      2873 => to_slv(opcode_type, 16#0A#),
      2874 => to_slv(opcode_type, 16#06#),
      2875 => to_slv(opcode_type, 16#0D#),
      2876 => to_slv(opcode_type, 16#0D#),
      2877 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#07#),
      2881 => to_slv(opcode_type, 16#06#),
      2882 => to_slv(opcode_type, 16#09#),
      2883 => to_slv(opcode_type, 16#08#),
      2884 => to_slv(opcode_type, 16#11#),
      2885 => to_slv(opcode_type, 16#21#),
      2886 => to_slv(opcode_type, 16#08#),
      2887 => to_slv(opcode_type, 16#0A#),
      2888 => to_slv(opcode_type, 16#0C#),
      2889 => to_slv(opcode_type, 16#08#),
      2890 => to_slv(opcode_type, 16#03#),
      2891 => to_slv(opcode_type, 16#94#),
      2892 => to_slv(opcode_type, 16#02#),
      2893 => to_slv(opcode_type, 16#11#),
      2894 => to_slv(opcode_type, 16#09#),
      2895 => to_slv(opcode_type, 16#08#),
      2896 => to_slv(opcode_type, 16#08#),
      2897 => to_slv(opcode_type, 16#0F#),
      2898 => to_slv(opcode_type, 16#11#),
      2899 => to_slv(opcode_type, 16#07#),
      2900 => to_slv(opcode_type, 16#0F#),
      2901 => to_slv(opcode_type, 16#0C#),
      2902 => to_slv(opcode_type, 16#08#),
      2903 => to_slv(opcode_type, 16#06#),
      2904 => to_slv(opcode_type, 16#0C#),
      2905 => to_slv(opcode_type, 16#0D#),
      2906 => to_slv(opcode_type, 16#07#),
      2907 => to_slv(opcode_type, 16#0D#),
      2908 => to_slv(opcode_type, 16#0C#),
      2909 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#08#),
      2913 => to_slv(opcode_type, 16#08#),
      2914 => to_slv(opcode_type, 16#06#),
      2915 => to_slv(opcode_type, 16#08#),
      2916 => to_slv(opcode_type, 16#0F#),
      2917 => to_slv(opcode_type, 16#0E#),
      2918 => to_slv(opcode_type, 16#09#),
      2919 => to_slv(opcode_type, 16#85#),
      2920 => to_slv(opcode_type, 16#11#),
      2921 => to_slv(opcode_type, 16#09#),
      2922 => to_slv(opcode_type, 16#07#),
      2923 => to_slv(opcode_type, 16#0A#),
      2924 => to_slv(opcode_type, 16#0A#),
      2925 => to_slv(opcode_type, 16#07#),
      2926 => to_slv(opcode_type, 16#10#),
      2927 => to_slv(opcode_type, 16#0F#),
      2928 => to_slv(opcode_type, 16#09#),
      2929 => to_slv(opcode_type, 16#07#),
      2930 => to_slv(opcode_type, 16#09#),
      2931 => to_slv(opcode_type, 16#0A#),
      2932 => to_slv(opcode_type, 16#0C#),
      2933 => to_slv(opcode_type, 16#08#),
      2934 => to_slv(opcode_type, 16#0C#),
      2935 => to_slv(opcode_type, 16#0D#),
      2936 => to_slv(opcode_type, 16#07#),
      2937 => to_slv(opcode_type, 16#09#),
      2938 => to_slv(opcode_type, 16#0F#),
      2939 => to_slv(opcode_type, 16#1C#),
      2940 => to_slv(opcode_type, 16#0F#),
      2941 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#09#),
      2945 => to_slv(opcode_type, 16#06#),
      2946 => to_slv(opcode_type, 16#06#),
      2947 => to_slv(opcode_type, 16#05#),
      2948 => to_slv(opcode_type, 16#0A#),
      2949 => to_slv(opcode_type, 16#08#),
      2950 => to_slv(opcode_type, 16#11#),
      2951 => to_slv(opcode_type, 16#0F#),
      2952 => to_slv(opcode_type, 16#08#),
      2953 => to_slv(opcode_type, 16#06#),
      2954 => to_slv(opcode_type, 16#0E#),
      2955 => to_slv(opcode_type, 16#0C#),
      2956 => to_slv(opcode_type, 16#02#),
      2957 => to_slv(opcode_type, 16#0B#),
      2958 => to_slv(opcode_type, 16#07#),
      2959 => to_slv(opcode_type, 16#09#),
      2960 => to_slv(opcode_type, 16#06#),
      2961 => to_slv(opcode_type, 16#0C#),
      2962 => to_slv(opcode_type, 16#0D#),
      2963 => to_slv(opcode_type, 16#08#),
      2964 => to_slv(opcode_type, 16#81#),
      2965 => to_slv(opcode_type, 16#0E#),
      2966 => to_slv(opcode_type, 16#08#),
      2967 => to_slv(opcode_type, 16#07#),
      2968 => to_slv(opcode_type, 16#0D#),
      2969 => to_slv(opcode_type, 16#0F#),
      2970 => to_slv(opcode_type, 16#09#),
      2971 => to_slv(opcode_type, 16#0C#),
      2972 => to_slv(opcode_type, 16#46#),
      2973 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#08#),
      2977 => to_slv(opcode_type, 16#08#),
      2978 => to_slv(opcode_type, 16#07#),
      2979 => to_slv(opcode_type, 16#01#),
      2980 => to_slv(opcode_type, 16#0D#),
      2981 => to_slv(opcode_type, 16#09#),
      2982 => to_slv(opcode_type, 16#0C#),
      2983 => to_slv(opcode_type, 16#10#),
      2984 => to_slv(opcode_type, 16#06#),
      2985 => to_slv(opcode_type, 16#07#),
      2986 => to_slv(opcode_type, 16#94#),
      2987 => to_slv(opcode_type, 16#0B#),
      2988 => to_slv(opcode_type, 16#09#),
      2989 => to_slv(opcode_type, 16#10#),
      2990 => to_slv(opcode_type, 16#0B#),
      2991 => to_slv(opcode_type, 16#09#),
      2992 => to_slv(opcode_type, 16#08#),
      2993 => to_slv(opcode_type, 16#03#),
      2994 => to_slv(opcode_type, 16#0F#),
      2995 => to_slv(opcode_type, 16#08#),
      2996 => to_slv(opcode_type, 16#0A#),
      2997 => to_slv(opcode_type, 16#0B#),
      2998 => to_slv(opcode_type, 16#06#),
      2999 => to_slv(opcode_type, 16#08#),
      3000 => to_slv(opcode_type, 16#0F#),
      3001 => to_slv(opcode_type, 16#0E#),
      3002 => to_slv(opcode_type, 16#06#),
      3003 => to_slv(opcode_type, 16#0A#),
      3004 => to_slv(opcode_type, 16#10#),
      3005 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#08#),
      3009 => to_slv(opcode_type, 16#07#),
      3010 => to_slv(opcode_type, 16#07#),
      3011 => to_slv(opcode_type, 16#01#),
      3012 => to_slv(opcode_type, 16#0C#),
      3013 => to_slv(opcode_type, 16#02#),
      3014 => to_slv(opcode_type, 16#0C#),
      3015 => to_slv(opcode_type, 16#07#),
      3016 => to_slv(opcode_type, 16#06#),
      3017 => to_slv(opcode_type, 16#AD#),
      3018 => to_slv(opcode_type, 16#0C#),
      3019 => to_slv(opcode_type, 16#06#),
      3020 => to_slv(opcode_type, 16#11#),
      3021 => to_slv(opcode_type, 16#0E#),
      3022 => to_slv(opcode_type, 16#07#),
      3023 => to_slv(opcode_type, 16#06#),
      3024 => to_slv(opcode_type, 16#07#),
      3025 => to_slv(opcode_type, 16#0C#),
      3026 => to_slv(opcode_type, 16#0B#),
      3027 => to_slv(opcode_type, 16#06#),
      3028 => to_slv(opcode_type, 16#0A#),
      3029 => to_slv(opcode_type, 16#0E#),
      3030 => to_slv(opcode_type, 16#08#),
      3031 => to_slv(opcode_type, 16#06#),
      3032 => to_slv(opcode_type, 16#0D#),
      3033 => to_slv(opcode_type, 16#0A#),
      3034 => to_slv(opcode_type, 16#09#),
      3035 => to_slv(opcode_type, 16#0C#),
      3036 => to_slv(opcode_type, 16#0B#),
      3037 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#07#),
      3041 => to_slv(opcode_type, 16#08#),
      3042 => to_slv(opcode_type, 16#09#),
      3043 => to_slv(opcode_type, 16#04#),
      3044 => to_slv(opcode_type, 16#0E#),
      3045 => to_slv(opcode_type, 16#06#),
      3046 => to_slv(opcode_type, 16#0B#),
      3047 => to_slv(opcode_type, 16#11#),
      3048 => to_slv(opcode_type, 16#08#),
      3049 => to_slv(opcode_type, 16#06#),
      3050 => to_slv(opcode_type, 16#11#),
      3051 => to_slv(opcode_type, 16#0B#),
      3052 => to_slv(opcode_type, 16#03#),
      3053 => to_slv(opcode_type, 16#0B#),
      3054 => to_slv(opcode_type, 16#06#),
      3055 => to_slv(opcode_type, 16#08#),
      3056 => to_slv(opcode_type, 16#08#),
      3057 => to_slv(opcode_type, 16#11#),
      3058 => to_slv(opcode_type, 16#7B#),
      3059 => to_slv(opcode_type, 16#09#),
      3060 => to_slv(opcode_type, 16#0B#),
      3061 => to_slv(opcode_type, 16#0D#),
      3062 => to_slv(opcode_type, 16#06#),
      3063 => to_slv(opcode_type, 16#07#),
      3064 => to_slv(opcode_type, 16#11#),
      3065 => to_slv(opcode_type, 16#0E#),
      3066 => to_slv(opcode_type, 16#09#),
      3067 => to_slv(opcode_type, 16#0C#),
      3068 => to_slv(opcode_type, 16#0C#),
      3069 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#08#),
      3073 => to_slv(opcode_type, 16#07#),
      3074 => to_slv(opcode_type, 16#06#),
      3075 => to_slv(opcode_type, 16#03#),
      3076 => to_slv(opcode_type, 16#0E#),
      3077 => to_slv(opcode_type, 16#07#),
      3078 => to_slv(opcode_type, 16#11#),
      3079 => to_slv(opcode_type, 16#CC#),
      3080 => to_slv(opcode_type, 16#06#),
      3081 => to_slv(opcode_type, 16#06#),
      3082 => to_slv(opcode_type, 16#0E#),
      3083 => to_slv(opcode_type, 16#0F#),
      3084 => to_slv(opcode_type, 16#05#),
      3085 => to_slv(opcode_type, 16#0B#),
      3086 => to_slv(opcode_type, 16#08#),
      3087 => to_slv(opcode_type, 16#06#),
      3088 => to_slv(opcode_type, 16#09#),
      3089 => to_slv(opcode_type, 16#10#),
      3090 => to_slv(opcode_type, 16#0B#),
      3091 => to_slv(opcode_type, 16#09#),
      3092 => to_slv(opcode_type, 16#0B#),
      3093 => to_slv(opcode_type, 16#0C#),
      3094 => to_slv(opcode_type, 16#06#),
      3095 => to_slv(opcode_type, 16#06#),
      3096 => to_slv(opcode_type, 16#0C#),
      3097 => to_slv(opcode_type, 16#0F#),
      3098 => to_slv(opcode_type, 16#06#),
      3099 => to_slv(opcode_type, 16#10#),
      3100 => to_slv(opcode_type, 16#EA#),
      3101 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#08#),
      3105 => to_slv(opcode_type, 16#08#),
      3106 => to_slv(opcode_type, 16#08#),
      3107 => to_slv(opcode_type, 16#06#),
      3108 => to_slv(opcode_type, 16#0F#),
      3109 => to_slv(opcode_type, 16#0E#),
      3110 => to_slv(opcode_type, 16#04#),
      3111 => to_slv(opcode_type, 16#0F#),
      3112 => to_slv(opcode_type, 16#09#),
      3113 => to_slv(opcode_type, 16#09#),
      3114 => to_slv(opcode_type, 16#0A#),
      3115 => to_slv(opcode_type, 16#10#),
      3116 => to_slv(opcode_type, 16#08#),
      3117 => to_slv(opcode_type, 16#0A#),
      3118 => to_slv(opcode_type, 16#0A#),
      3119 => to_slv(opcode_type, 16#06#),
      3120 => to_slv(opcode_type, 16#09#),
      3121 => to_slv(opcode_type, 16#03#),
      3122 => to_slv(opcode_type, 16#0E#),
      3123 => to_slv(opcode_type, 16#07#),
      3124 => to_slv(opcode_type, 16#87#),
      3125 => to_slv(opcode_type, 16#0A#),
      3126 => to_slv(opcode_type, 16#09#),
      3127 => to_slv(opcode_type, 16#08#),
      3128 => to_slv(opcode_type, 16#0F#),
      3129 => to_slv(opcode_type, 16#10#),
      3130 => to_slv(opcode_type, 16#07#),
      3131 => to_slv(opcode_type, 16#7D#),
      3132 => to_slv(opcode_type, 16#0E#),
      3133 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#06#),
      3137 => to_slv(opcode_type, 16#08#),
      3138 => to_slv(opcode_type, 16#08#),
      3139 => to_slv(opcode_type, 16#06#),
      3140 => to_slv(opcode_type, 16#0C#),
      3141 => to_slv(opcode_type, 16#0B#),
      3142 => to_slv(opcode_type, 16#05#),
      3143 => to_slv(opcode_type, 16#0C#),
      3144 => to_slv(opcode_type, 16#09#),
      3145 => to_slv(opcode_type, 16#08#),
      3146 => to_slv(opcode_type, 16#11#),
      3147 => to_slv(opcode_type, 16#10#),
      3148 => to_slv(opcode_type, 16#09#),
      3149 => to_slv(opcode_type, 16#0A#),
      3150 => to_slv(opcode_type, 16#0F#),
      3151 => to_slv(opcode_type, 16#06#),
      3152 => to_slv(opcode_type, 16#07#),
      3153 => to_slv(opcode_type, 16#03#),
      3154 => to_slv(opcode_type, 16#11#),
      3155 => to_slv(opcode_type, 16#08#),
      3156 => to_slv(opcode_type, 16#0A#),
      3157 => to_slv(opcode_type, 16#0F#),
      3158 => to_slv(opcode_type, 16#09#),
      3159 => to_slv(opcode_type, 16#09#),
      3160 => to_slv(opcode_type, 16#0F#),
      3161 => to_slv(opcode_type, 16#11#),
      3162 => to_slv(opcode_type, 16#09#),
      3163 => to_slv(opcode_type, 16#0D#),
      3164 => to_slv(opcode_type, 16#0D#),
      3165 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#09#),
      3169 => to_slv(opcode_type, 16#07#),
      3170 => to_slv(opcode_type, 16#08#),
      3171 => to_slv(opcode_type, 16#05#),
      3172 => to_slv(opcode_type, 16#0C#),
      3173 => to_slv(opcode_type, 16#05#),
      3174 => to_slv(opcode_type, 16#0D#),
      3175 => to_slv(opcode_type, 16#09#),
      3176 => to_slv(opcode_type, 16#09#),
      3177 => to_slv(opcode_type, 16#0C#),
      3178 => to_slv(opcode_type, 16#0B#),
      3179 => to_slv(opcode_type, 16#08#),
      3180 => to_slv(opcode_type, 16#0E#),
      3181 => to_slv(opcode_type, 16#0E#),
      3182 => to_slv(opcode_type, 16#09#),
      3183 => to_slv(opcode_type, 16#08#),
      3184 => to_slv(opcode_type, 16#07#),
      3185 => to_slv(opcode_type, 16#0F#),
      3186 => to_slv(opcode_type, 16#0A#),
      3187 => to_slv(opcode_type, 16#06#),
      3188 => to_slv(opcode_type, 16#11#),
      3189 => to_slv(opcode_type, 16#11#),
      3190 => to_slv(opcode_type, 16#07#),
      3191 => to_slv(opcode_type, 16#09#),
      3192 => to_slv(opcode_type, 16#10#),
      3193 => to_slv(opcode_type, 16#0E#),
      3194 => to_slv(opcode_type, 16#08#),
      3195 => to_slv(opcode_type, 16#0D#),
      3196 => to_slv(opcode_type, 16#0D#),
      3197 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#08#),
      3201 => to_slv(opcode_type, 16#08#),
      3202 => to_slv(opcode_type, 16#06#),
      3203 => to_slv(opcode_type, 16#06#),
      3204 => to_slv(opcode_type, 16#11#),
      3205 => to_slv(opcode_type, 16#0E#),
      3206 => to_slv(opcode_type, 16#07#),
      3207 => to_slv(opcode_type, 16#0A#),
      3208 => to_slv(opcode_type, 16#0A#),
      3209 => to_slv(opcode_type, 16#07#),
      3210 => to_slv(opcode_type, 16#03#),
      3211 => to_slv(opcode_type, 16#0D#),
      3212 => to_slv(opcode_type, 16#01#),
      3213 => to_slv(opcode_type, 16#11#),
      3214 => to_slv(opcode_type, 16#06#),
      3215 => to_slv(opcode_type, 16#08#),
      3216 => to_slv(opcode_type, 16#06#),
      3217 => to_slv(opcode_type, 16#0C#),
      3218 => to_slv(opcode_type, 16#2D#),
      3219 => to_slv(opcode_type, 16#09#),
      3220 => to_slv(opcode_type, 16#0C#),
      3221 => to_slv(opcode_type, 16#11#),
      3222 => to_slv(opcode_type, 16#06#),
      3223 => to_slv(opcode_type, 16#07#),
      3224 => to_slv(opcode_type, 16#0D#),
      3225 => to_slv(opcode_type, 16#0D#),
      3226 => to_slv(opcode_type, 16#06#),
      3227 => to_slv(opcode_type, 16#6C#),
      3228 => to_slv(opcode_type, 16#0E#),
      3229 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#09#),
      3234 => to_slv(opcode_type, 16#06#),
      3235 => to_slv(opcode_type, 16#02#),
      3236 => to_slv(opcode_type, 16#0A#),
      3237 => to_slv(opcode_type, 16#03#),
      3238 => to_slv(opcode_type, 16#0F#),
      3239 => to_slv(opcode_type, 16#07#),
      3240 => to_slv(opcode_type, 16#09#),
      3241 => to_slv(opcode_type, 16#10#),
      3242 => to_slv(opcode_type, 16#0B#),
      3243 => to_slv(opcode_type, 16#07#),
      3244 => to_slv(opcode_type, 16#0E#),
      3245 => to_slv(opcode_type, 16#0D#),
      3246 => to_slv(opcode_type, 16#07#),
      3247 => to_slv(opcode_type, 16#09#),
      3248 => to_slv(opcode_type, 16#06#),
      3249 => to_slv(opcode_type, 16#5A#),
      3250 => to_slv(opcode_type, 16#0F#),
      3251 => to_slv(opcode_type, 16#09#),
      3252 => to_slv(opcode_type, 16#0E#),
      3253 => to_slv(opcode_type, 16#0A#),
      3254 => to_slv(opcode_type, 16#08#),
      3255 => to_slv(opcode_type, 16#07#),
      3256 => to_slv(opcode_type, 16#0C#),
      3257 => to_slv(opcode_type, 16#11#),
      3258 => to_slv(opcode_type, 16#08#),
      3259 => to_slv(opcode_type, 16#0D#),
      3260 => to_slv(opcode_type, 16#0F#),
      3261 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#08#),
      3265 => to_slv(opcode_type, 16#07#),
      3266 => to_slv(opcode_type, 16#07#),
      3267 => to_slv(opcode_type, 16#05#),
      3268 => to_slv(opcode_type, 16#11#),
      3269 => to_slv(opcode_type, 16#06#),
      3270 => to_slv(opcode_type, 16#0F#),
      3271 => to_slv(opcode_type, 16#EE#),
      3272 => to_slv(opcode_type, 16#06#),
      3273 => to_slv(opcode_type, 16#09#),
      3274 => to_slv(opcode_type, 16#0D#),
      3275 => to_slv(opcode_type, 16#11#),
      3276 => to_slv(opcode_type, 16#06#),
      3277 => to_slv(opcode_type, 16#0B#),
      3278 => to_slv(opcode_type, 16#BA#),
      3279 => to_slv(opcode_type, 16#09#),
      3280 => to_slv(opcode_type, 16#09#),
      3281 => to_slv(opcode_type, 16#05#),
      3282 => to_slv(opcode_type, 16#42#),
      3283 => to_slv(opcode_type, 16#09#),
      3284 => to_slv(opcode_type, 16#0A#),
      3285 => to_slv(opcode_type, 16#0F#),
      3286 => to_slv(opcode_type, 16#06#),
      3287 => to_slv(opcode_type, 16#07#),
      3288 => to_slv(opcode_type, 16#0D#),
      3289 => to_slv(opcode_type, 16#0E#),
      3290 => to_slv(opcode_type, 16#06#),
      3291 => to_slv(opcode_type, 16#10#),
      3292 => to_slv(opcode_type, 16#0A#),
      3293 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#06#),
      3297 => to_slv(opcode_type, 16#08#),
      3298 => to_slv(opcode_type, 16#08#),
      3299 => to_slv(opcode_type, 16#06#),
      3300 => to_slv(opcode_type, 16#10#),
      3301 => to_slv(opcode_type, 16#11#),
      3302 => to_slv(opcode_type, 16#02#),
      3303 => to_slv(opcode_type, 16#0E#),
      3304 => to_slv(opcode_type, 16#08#),
      3305 => to_slv(opcode_type, 16#03#),
      3306 => to_slv(opcode_type, 16#0B#),
      3307 => to_slv(opcode_type, 16#09#),
      3308 => to_slv(opcode_type, 16#10#),
      3309 => to_slv(opcode_type, 16#0A#),
      3310 => to_slv(opcode_type, 16#09#),
      3311 => to_slv(opcode_type, 16#09#),
      3312 => to_slv(opcode_type, 16#07#),
      3313 => to_slv(opcode_type, 16#F8#),
      3314 => to_slv(opcode_type, 16#0E#),
      3315 => to_slv(opcode_type, 16#09#),
      3316 => to_slv(opcode_type, 16#11#),
      3317 => to_slv(opcode_type, 16#0D#),
      3318 => to_slv(opcode_type, 16#06#),
      3319 => to_slv(opcode_type, 16#07#),
      3320 => to_slv(opcode_type, 16#0B#),
      3321 => to_slv(opcode_type, 16#28#),
      3322 => to_slv(opcode_type, 16#07#),
      3323 => to_slv(opcode_type, 16#10#),
      3324 => to_slv(opcode_type, 16#0E#),
      3325 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#06#),
      3329 => to_slv(opcode_type, 16#06#),
      3330 => to_slv(opcode_type, 16#09#),
      3331 => to_slv(opcode_type, 16#07#),
      3332 => to_slv(opcode_type, 16#0E#),
      3333 => to_slv(opcode_type, 16#0A#),
      3334 => to_slv(opcode_type, 16#07#),
      3335 => to_slv(opcode_type, 16#0D#),
      3336 => to_slv(opcode_type, 16#0D#),
      3337 => to_slv(opcode_type, 16#09#),
      3338 => to_slv(opcode_type, 16#08#),
      3339 => to_slv(opcode_type, 16#AF#),
      3340 => to_slv(opcode_type, 16#10#),
      3341 => to_slv(opcode_type, 16#08#),
      3342 => to_slv(opcode_type, 16#11#),
      3343 => to_slv(opcode_type, 16#0F#),
      3344 => to_slv(opcode_type, 16#07#),
      3345 => to_slv(opcode_type, 16#09#),
      3346 => to_slv(opcode_type, 16#06#),
      3347 => to_slv(opcode_type, 16#0E#),
      3348 => to_slv(opcode_type, 16#0D#),
      3349 => to_slv(opcode_type, 16#06#),
      3350 => to_slv(opcode_type, 16#0C#),
      3351 => to_slv(opcode_type, 16#0A#),
      3352 => to_slv(opcode_type, 16#06#),
      3353 => to_slv(opcode_type, 16#07#),
      3354 => to_slv(opcode_type, 16#10#),
      3355 => to_slv(opcode_type, 16#10#),
      3356 => to_slv(opcode_type, 16#10#),
      3357 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#07#),
      3361 => to_slv(opcode_type, 16#09#),
      3362 => to_slv(opcode_type, 16#09#),
      3363 => to_slv(opcode_type, 16#01#),
      3364 => to_slv(opcode_type, 16#0D#),
      3365 => to_slv(opcode_type, 16#09#),
      3366 => to_slv(opcode_type, 16#0F#),
      3367 => to_slv(opcode_type, 16#41#),
      3368 => to_slv(opcode_type, 16#07#),
      3369 => to_slv(opcode_type, 16#07#),
      3370 => to_slv(opcode_type, 16#0B#),
      3371 => to_slv(opcode_type, 16#0D#),
      3372 => to_slv(opcode_type, 16#07#),
      3373 => to_slv(opcode_type, 16#0C#),
      3374 => to_slv(opcode_type, 16#0E#),
      3375 => to_slv(opcode_type, 16#08#),
      3376 => to_slv(opcode_type, 16#08#),
      3377 => to_slv(opcode_type, 16#09#),
      3378 => to_slv(opcode_type, 16#0E#),
      3379 => to_slv(opcode_type, 16#0D#),
      3380 => to_slv(opcode_type, 16#06#),
      3381 => to_slv(opcode_type, 16#11#),
      3382 => to_slv(opcode_type, 16#0D#),
      3383 => to_slv(opcode_type, 16#09#),
      3384 => to_slv(opcode_type, 16#03#),
      3385 => to_slv(opcode_type, 16#0B#),
      3386 => to_slv(opcode_type, 16#07#),
      3387 => to_slv(opcode_type, 16#0E#),
      3388 => to_slv(opcode_type, 16#73#),
      3389 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#08#),
      3393 => to_slv(opcode_type, 16#09#),
      3394 => to_slv(opcode_type, 16#07#),
      3395 => to_slv(opcode_type, 16#03#),
      3396 => to_slv(opcode_type, 16#0A#),
      3397 => to_slv(opcode_type, 16#03#),
      3398 => to_slv(opcode_type, 16#0A#),
      3399 => to_slv(opcode_type, 16#08#),
      3400 => to_slv(opcode_type, 16#09#),
      3401 => to_slv(opcode_type, 16#0C#),
      3402 => to_slv(opcode_type, 16#0C#),
      3403 => to_slv(opcode_type, 16#07#),
      3404 => to_slv(opcode_type, 16#0D#),
      3405 => to_slv(opcode_type, 16#0A#),
      3406 => to_slv(opcode_type, 16#06#),
      3407 => to_slv(opcode_type, 16#06#),
      3408 => to_slv(opcode_type, 16#07#),
      3409 => to_slv(opcode_type, 16#0E#),
      3410 => to_slv(opcode_type, 16#11#),
      3411 => to_slv(opcode_type, 16#08#),
      3412 => to_slv(opcode_type, 16#10#),
      3413 => to_slv(opcode_type, 16#11#),
      3414 => to_slv(opcode_type, 16#07#),
      3415 => to_slv(opcode_type, 16#08#),
      3416 => to_slv(opcode_type, 16#0A#),
      3417 => to_slv(opcode_type, 16#0F#),
      3418 => to_slv(opcode_type, 16#06#),
      3419 => to_slv(opcode_type, 16#0C#),
      3420 => to_slv(opcode_type, 16#0B#),
      3421 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#07#),
      3425 => to_slv(opcode_type, 16#06#),
      3426 => to_slv(opcode_type, 16#08#),
      3427 => to_slv(opcode_type, 16#02#),
      3428 => to_slv(opcode_type, 16#0B#),
      3429 => to_slv(opcode_type, 16#05#),
      3430 => to_slv(opcode_type, 16#11#),
      3431 => to_slv(opcode_type, 16#06#),
      3432 => to_slv(opcode_type, 16#06#),
      3433 => to_slv(opcode_type, 16#0B#),
      3434 => to_slv(opcode_type, 16#0A#),
      3435 => to_slv(opcode_type, 16#08#),
      3436 => to_slv(opcode_type, 16#0E#),
      3437 => to_slv(opcode_type, 16#10#),
      3438 => to_slv(opcode_type, 16#08#),
      3439 => to_slv(opcode_type, 16#07#),
      3440 => to_slv(opcode_type, 16#07#),
      3441 => to_slv(opcode_type, 16#0F#),
      3442 => to_slv(opcode_type, 16#11#),
      3443 => to_slv(opcode_type, 16#08#),
      3444 => to_slv(opcode_type, 16#0E#),
      3445 => to_slv(opcode_type, 16#0E#),
      3446 => to_slv(opcode_type, 16#06#),
      3447 => to_slv(opcode_type, 16#09#),
      3448 => to_slv(opcode_type, 16#0B#),
      3449 => to_slv(opcode_type, 16#22#),
      3450 => to_slv(opcode_type, 16#07#),
      3451 => to_slv(opcode_type, 16#10#),
      3452 => to_slv(opcode_type, 16#0A#),
      3453 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#08#),
      3457 => to_slv(opcode_type, 16#06#),
      3458 => to_slv(opcode_type, 16#08#),
      3459 => to_slv(opcode_type, 16#07#),
      3460 => to_slv(opcode_type, 16#0E#),
      3461 => to_slv(opcode_type, 16#11#),
      3462 => to_slv(opcode_type, 16#01#),
      3463 => to_slv(opcode_type, 16#0E#),
      3464 => to_slv(opcode_type, 16#06#),
      3465 => to_slv(opcode_type, 16#04#),
      3466 => to_slv(opcode_type, 16#EB#),
      3467 => to_slv(opcode_type, 16#07#),
      3468 => to_slv(opcode_type, 16#0C#),
      3469 => to_slv(opcode_type, 16#11#),
      3470 => to_slv(opcode_type, 16#08#),
      3471 => to_slv(opcode_type, 16#06#),
      3472 => to_slv(opcode_type, 16#08#),
      3473 => to_slv(opcode_type, 16#0A#),
      3474 => to_slv(opcode_type, 16#0D#),
      3475 => to_slv(opcode_type, 16#06#),
      3476 => to_slv(opcode_type, 16#0F#),
      3477 => to_slv(opcode_type, 16#0C#),
      3478 => to_slv(opcode_type, 16#06#),
      3479 => to_slv(opcode_type, 16#08#),
      3480 => to_slv(opcode_type, 16#0C#),
      3481 => to_slv(opcode_type, 16#10#),
      3482 => to_slv(opcode_type, 16#08#),
      3483 => to_slv(opcode_type, 16#0F#),
      3484 => to_slv(opcode_type, 16#0A#),
      3485 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#06#),
      3489 => to_slv(opcode_type, 16#08#),
      3490 => to_slv(opcode_type, 16#06#),
      3491 => to_slv(opcode_type, 16#01#),
      3492 => to_slv(opcode_type, 16#0F#),
      3493 => to_slv(opcode_type, 16#06#),
      3494 => to_slv(opcode_type, 16#0A#),
      3495 => to_slv(opcode_type, 16#11#),
      3496 => to_slv(opcode_type, 16#09#),
      3497 => to_slv(opcode_type, 16#07#),
      3498 => to_slv(opcode_type, 16#0E#),
      3499 => to_slv(opcode_type, 16#0A#),
      3500 => to_slv(opcode_type, 16#07#),
      3501 => to_slv(opcode_type, 16#0F#),
      3502 => to_slv(opcode_type, 16#0E#),
      3503 => to_slv(opcode_type, 16#08#),
      3504 => to_slv(opcode_type, 16#06#),
      3505 => to_slv(opcode_type, 16#04#),
      3506 => to_slv(opcode_type, 16#F1#),
      3507 => to_slv(opcode_type, 16#06#),
      3508 => to_slv(opcode_type, 16#44#),
      3509 => to_slv(opcode_type, 16#0B#),
      3510 => to_slv(opcode_type, 16#08#),
      3511 => to_slv(opcode_type, 16#06#),
      3512 => to_slv(opcode_type, 16#11#),
      3513 => to_slv(opcode_type, 16#0A#),
      3514 => to_slv(opcode_type, 16#09#),
      3515 => to_slv(opcode_type, 16#0C#),
      3516 => to_slv(opcode_type, 16#0C#),
      3517 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#06#),
      3521 => to_slv(opcode_type, 16#08#),
      3522 => to_slv(opcode_type, 16#07#),
      3523 => to_slv(opcode_type, 16#08#),
      3524 => to_slv(opcode_type, 16#0A#),
      3525 => to_slv(opcode_type, 16#0E#),
      3526 => to_slv(opcode_type, 16#03#),
      3527 => to_slv(opcode_type, 16#3F#),
      3528 => to_slv(opcode_type, 16#07#),
      3529 => to_slv(opcode_type, 16#06#),
      3530 => to_slv(opcode_type, 16#0C#),
      3531 => to_slv(opcode_type, 16#0F#),
      3532 => to_slv(opcode_type, 16#04#),
      3533 => to_slv(opcode_type, 16#0D#),
      3534 => to_slv(opcode_type, 16#07#),
      3535 => to_slv(opcode_type, 16#07#),
      3536 => to_slv(opcode_type, 16#06#),
      3537 => to_slv(opcode_type, 16#0D#),
      3538 => to_slv(opcode_type, 16#0F#),
      3539 => to_slv(opcode_type, 16#07#),
      3540 => to_slv(opcode_type, 16#0D#),
      3541 => to_slv(opcode_type, 16#0A#),
      3542 => to_slv(opcode_type, 16#08#),
      3543 => to_slv(opcode_type, 16#08#),
      3544 => to_slv(opcode_type, 16#0A#),
      3545 => to_slv(opcode_type, 16#10#),
      3546 => to_slv(opcode_type, 16#09#),
      3547 => to_slv(opcode_type, 16#0C#),
      3548 => to_slv(opcode_type, 16#0D#),
      3549 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#09#),
      3553 => to_slv(opcode_type, 16#08#),
      3554 => to_slv(opcode_type, 16#08#),
      3555 => to_slv(opcode_type, 16#02#),
      3556 => to_slv(opcode_type, 16#0F#),
      3557 => to_slv(opcode_type, 16#09#),
      3558 => to_slv(opcode_type, 16#0B#),
      3559 => to_slv(opcode_type, 16#0C#),
      3560 => to_slv(opcode_type, 16#06#),
      3561 => to_slv(opcode_type, 16#08#),
      3562 => to_slv(opcode_type, 16#11#),
      3563 => to_slv(opcode_type, 16#0E#),
      3564 => to_slv(opcode_type, 16#04#),
      3565 => to_slv(opcode_type, 16#0F#),
      3566 => to_slv(opcode_type, 16#09#),
      3567 => to_slv(opcode_type, 16#07#),
      3568 => to_slv(opcode_type, 16#09#),
      3569 => to_slv(opcode_type, 16#10#),
      3570 => to_slv(opcode_type, 16#0F#),
      3571 => to_slv(opcode_type, 16#06#),
      3572 => to_slv(opcode_type, 16#0E#),
      3573 => to_slv(opcode_type, 16#0F#),
      3574 => to_slv(opcode_type, 16#06#),
      3575 => to_slv(opcode_type, 16#06#),
      3576 => to_slv(opcode_type, 16#0D#),
      3577 => to_slv(opcode_type, 16#11#),
      3578 => to_slv(opcode_type, 16#09#),
      3579 => to_slv(opcode_type, 16#0E#),
      3580 => to_slv(opcode_type, 16#0C#),
      3581 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#09#),
      3585 => to_slv(opcode_type, 16#06#),
      3586 => to_slv(opcode_type, 16#07#),
      3587 => to_slv(opcode_type, 16#09#),
      3588 => to_slv(opcode_type, 16#0C#),
      3589 => to_slv(opcode_type, 16#72#),
      3590 => to_slv(opcode_type, 16#09#),
      3591 => to_slv(opcode_type, 16#10#),
      3592 => to_slv(opcode_type, 16#0A#),
      3593 => to_slv(opcode_type, 16#09#),
      3594 => to_slv(opcode_type, 16#05#),
      3595 => to_slv(opcode_type, 16#0D#),
      3596 => to_slv(opcode_type, 16#02#),
      3597 => to_slv(opcode_type, 16#0B#),
      3598 => to_slv(opcode_type, 16#06#),
      3599 => to_slv(opcode_type, 16#07#),
      3600 => to_slv(opcode_type, 16#06#),
      3601 => to_slv(opcode_type, 16#0D#),
      3602 => to_slv(opcode_type, 16#51#),
      3603 => to_slv(opcode_type, 16#06#),
      3604 => to_slv(opcode_type, 16#0B#),
      3605 => to_slv(opcode_type, 16#0E#),
      3606 => to_slv(opcode_type, 16#06#),
      3607 => to_slv(opcode_type, 16#09#),
      3608 => to_slv(opcode_type, 16#0D#),
      3609 => to_slv(opcode_type, 16#0E#),
      3610 => to_slv(opcode_type, 16#06#),
      3611 => to_slv(opcode_type, 16#5E#),
      3612 => to_slv(opcode_type, 16#0E#),
      3613 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#06#),
      3617 => to_slv(opcode_type, 16#09#),
      3618 => to_slv(opcode_type, 16#09#),
      3619 => to_slv(opcode_type, 16#01#),
      3620 => to_slv(opcode_type, 16#0E#),
      3621 => to_slv(opcode_type, 16#05#),
      3622 => to_slv(opcode_type, 16#0F#),
      3623 => to_slv(opcode_type, 16#08#),
      3624 => to_slv(opcode_type, 16#08#),
      3625 => to_slv(opcode_type, 16#48#),
      3626 => to_slv(opcode_type, 16#0A#),
      3627 => to_slv(opcode_type, 16#09#),
      3628 => to_slv(opcode_type, 16#11#),
      3629 => to_slv(opcode_type, 16#11#),
      3630 => to_slv(opcode_type, 16#09#),
      3631 => to_slv(opcode_type, 16#09#),
      3632 => to_slv(opcode_type, 16#09#),
      3633 => to_slv(opcode_type, 16#11#),
      3634 => to_slv(opcode_type, 16#1B#),
      3635 => to_slv(opcode_type, 16#07#),
      3636 => to_slv(opcode_type, 16#10#),
      3637 => to_slv(opcode_type, 16#0B#),
      3638 => to_slv(opcode_type, 16#09#),
      3639 => to_slv(opcode_type, 16#09#),
      3640 => to_slv(opcode_type, 16#0A#),
      3641 => to_slv(opcode_type, 16#0C#),
      3642 => to_slv(opcode_type, 16#08#),
      3643 => to_slv(opcode_type, 16#11#),
      3644 => to_slv(opcode_type, 16#0C#),
      3645 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#06#),
      3649 => to_slv(opcode_type, 16#07#),
      3650 => to_slv(opcode_type, 16#07#),
      3651 => to_slv(opcode_type, 16#01#),
      3652 => to_slv(opcode_type, 16#0A#),
      3653 => to_slv(opcode_type, 16#04#),
      3654 => to_slv(opcode_type, 16#0A#),
      3655 => to_slv(opcode_type, 16#06#),
      3656 => to_slv(opcode_type, 16#06#),
      3657 => to_slv(opcode_type, 16#0D#),
      3658 => to_slv(opcode_type, 16#11#),
      3659 => to_slv(opcode_type, 16#09#),
      3660 => to_slv(opcode_type, 16#0B#),
      3661 => to_slv(opcode_type, 16#4B#),
      3662 => to_slv(opcode_type, 16#08#),
      3663 => to_slv(opcode_type, 16#08#),
      3664 => to_slv(opcode_type, 16#07#),
      3665 => to_slv(opcode_type, 16#11#),
      3666 => to_slv(opcode_type, 16#D2#),
      3667 => to_slv(opcode_type, 16#06#),
      3668 => to_slv(opcode_type, 16#10#),
      3669 => to_slv(opcode_type, 16#0C#),
      3670 => to_slv(opcode_type, 16#07#),
      3671 => to_slv(opcode_type, 16#09#),
      3672 => to_slv(opcode_type, 16#81#),
      3673 => to_slv(opcode_type, 16#0D#),
      3674 => to_slv(opcode_type, 16#09#),
      3675 => to_slv(opcode_type, 16#0A#),
      3676 => to_slv(opcode_type, 16#0B#),
      3677 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#07#),
      3681 => to_slv(opcode_type, 16#08#),
      3682 => to_slv(opcode_type, 16#07#),
      3683 => to_slv(opcode_type, 16#01#),
      3684 => to_slv(opcode_type, 16#0D#),
      3685 => to_slv(opcode_type, 16#04#),
      3686 => to_slv(opcode_type, 16#B4#),
      3687 => to_slv(opcode_type, 16#08#),
      3688 => to_slv(opcode_type, 16#06#),
      3689 => to_slv(opcode_type, 16#0B#),
      3690 => to_slv(opcode_type, 16#0B#),
      3691 => to_slv(opcode_type, 16#08#),
      3692 => to_slv(opcode_type, 16#0C#),
      3693 => to_slv(opcode_type, 16#0B#),
      3694 => to_slv(opcode_type, 16#07#),
      3695 => to_slv(opcode_type, 16#09#),
      3696 => to_slv(opcode_type, 16#06#),
      3697 => to_slv(opcode_type, 16#0A#),
      3698 => to_slv(opcode_type, 16#0B#),
      3699 => to_slv(opcode_type, 16#09#),
      3700 => to_slv(opcode_type, 16#0B#),
      3701 => to_slv(opcode_type, 16#0D#),
      3702 => to_slv(opcode_type, 16#08#),
      3703 => to_slv(opcode_type, 16#08#),
      3704 => to_slv(opcode_type, 16#10#),
      3705 => to_slv(opcode_type, 16#0A#),
      3706 => to_slv(opcode_type, 16#07#),
      3707 => to_slv(opcode_type, 16#0D#),
      3708 => to_slv(opcode_type, 16#0A#),
      3709 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#08#),
      3713 => to_slv(opcode_type, 16#09#),
      3714 => to_slv(opcode_type, 16#09#),
      3715 => to_slv(opcode_type, 16#04#),
      3716 => to_slv(opcode_type, 16#0A#),
      3717 => to_slv(opcode_type, 16#05#),
      3718 => to_slv(opcode_type, 16#9A#),
      3719 => to_slv(opcode_type, 16#08#),
      3720 => to_slv(opcode_type, 16#09#),
      3721 => to_slv(opcode_type, 16#0D#),
      3722 => to_slv(opcode_type, 16#11#),
      3723 => to_slv(opcode_type, 16#06#),
      3724 => to_slv(opcode_type, 16#0A#),
      3725 => to_slv(opcode_type, 16#0D#),
      3726 => to_slv(opcode_type, 16#08#),
      3727 => to_slv(opcode_type, 16#09#),
      3728 => to_slv(opcode_type, 16#08#),
      3729 => to_slv(opcode_type, 16#0D#),
      3730 => to_slv(opcode_type, 16#0A#),
      3731 => to_slv(opcode_type, 16#07#),
      3732 => to_slv(opcode_type, 16#0D#),
      3733 => to_slv(opcode_type, 16#0C#),
      3734 => to_slv(opcode_type, 16#06#),
      3735 => to_slv(opcode_type, 16#06#),
      3736 => to_slv(opcode_type, 16#10#),
      3737 => to_slv(opcode_type, 16#11#),
      3738 => to_slv(opcode_type, 16#08#),
      3739 => to_slv(opcode_type, 16#0B#),
      3740 => to_slv(opcode_type, 16#6E#),
      3741 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#06#),
      3745 => to_slv(opcode_type, 16#09#),
      3746 => to_slv(opcode_type, 16#09#),
      3747 => to_slv(opcode_type, 16#02#),
      3748 => to_slv(opcode_type, 16#0C#),
      3749 => to_slv(opcode_type, 16#08#),
      3750 => to_slv(opcode_type, 16#0B#),
      3751 => to_slv(opcode_type, 16#0C#),
      3752 => to_slv(opcode_type, 16#07#),
      3753 => to_slv(opcode_type, 16#03#),
      3754 => to_slv(opcode_type, 16#2C#),
      3755 => to_slv(opcode_type, 16#08#),
      3756 => to_slv(opcode_type, 16#0E#),
      3757 => to_slv(opcode_type, 16#11#),
      3758 => to_slv(opcode_type, 16#07#),
      3759 => to_slv(opcode_type, 16#06#),
      3760 => to_slv(opcode_type, 16#06#),
      3761 => to_slv(opcode_type, 16#0D#),
      3762 => to_slv(opcode_type, 16#11#),
      3763 => to_slv(opcode_type, 16#08#),
      3764 => to_slv(opcode_type, 16#0B#),
      3765 => to_slv(opcode_type, 16#0F#),
      3766 => to_slv(opcode_type, 16#09#),
      3767 => to_slv(opcode_type, 16#09#),
      3768 => to_slv(opcode_type, 16#27#),
      3769 => to_slv(opcode_type, 16#82#),
      3770 => to_slv(opcode_type, 16#09#),
      3771 => to_slv(opcode_type, 16#0A#),
      3772 => to_slv(opcode_type, 16#0B#),
      3773 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#07#),
      3777 => to_slv(opcode_type, 16#09#),
      3778 => to_slv(opcode_type, 16#08#),
      3779 => to_slv(opcode_type, 16#04#),
      3780 => to_slv(opcode_type, 16#0C#),
      3781 => to_slv(opcode_type, 16#02#),
      3782 => to_slv(opcode_type, 16#0E#),
      3783 => to_slv(opcode_type, 16#08#),
      3784 => to_slv(opcode_type, 16#07#),
      3785 => to_slv(opcode_type, 16#0E#),
      3786 => to_slv(opcode_type, 16#10#),
      3787 => to_slv(opcode_type, 16#06#),
      3788 => to_slv(opcode_type, 16#11#),
      3789 => to_slv(opcode_type, 16#0F#),
      3790 => to_slv(opcode_type, 16#08#),
      3791 => to_slv(opcode_type, 16#06#),
      3792 => to_slv(opcode_type, 16#07#),
      3793 => to_slv(opcode_type, 16#0F#),
      3794 => to_slv(opcode_type, 16#0A#),
      3795 => to_slv(opcode_type, 16#06#),
      3796 => to_slv(opcode_type, 16#0E#),
      3797 => to_slv(opcode_type, 16#0D#),
      3798 => to_slv(opcode_type, 16#07#),
      3799 => to_slv(opcode_type, 16#08#),
      3800 => to_slv(opcode_type, 16#10#),
      3801 => to_slv(opcode_type, 16#10#),
      3802 => to_slv(opcode_type, 16#06#),
      3803 => to_slv(opcode_type, 16#10#),
      3804 => to_slv(opcode_type, 16#0E#),
      3805 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#09#),
      3809 => to_slv(opcode_type, 16#07#),
      3810 => to_slv(opcode_type, 16#06#),
      3811 => to_slv(opcode_type, 16#02#),
      3812 => to_slv(opcode_type, 16#0C#),
      3813 => to_slv(opcode_type, 16#05#),
      3814 => to_slv(opcode_type, 16#0F#),
      3815 => to_slv(opcode_type, 16#09#),
      3816 => to_slv(opcode_type, 16#06#),
      3817 => to_slv(opcode_type, 16#3A#),
      3818 => to_slv(opcode_type, 16#10#),
      3819 => to_slv(opcode_type, 16#06#),
      3820 => to_slv(opcode_type, 16#0B#),
      3821 => to_slv(opcode_type, 16#0B#),
      3822 => to_slv(opcode_type, 16#09#),
      3823 => to_slv(opcode_type, 16#09#),
      3824 => to_slv(opcode_type, 16#08#),
      3825 => to_slv(opcode_type, 16#0B#),
      3826 => to_slv(opcode_type, 16#0D#),
      3827 => to_slv(opcode_type, 16#09#),
      3828 => to_slv(opcode_type, 16#0F#),
      3829 => to_slv(opcode_type, 16#B0#),
      3830 => to_slv(opcode_type, 16#09#),
      3831 => to_slv(opcode_type, 16#07#),
      3832 => to_slv(opcode_type, 16#10#),
      3833 => to_slv(opcode_type, 16#0E#),
      3834 => to_slv(opcode_type, 16#07#),
      3835 => to_slv(opcode_type, 16#10#),
      3836 => to_slv(opcode_type, 16#72#),
      3837 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#06#),
      3841 => to_slv(opcode_type, 16#07#),
      3842 => to_slv(opcode_type, 16#07#),
      3843 => to_slv(opcode_type, 16#09#),
      3844 => to_slv(opcode_type, 16#10#),
      3845 => to_slv(opcode_type, 16#0E#),
      3846 => to_slv(opcode_type, 16#01#),
      3847 => to_slv(opcode_type, 16#0A#),
      3848 => to_slv(opcode_type, 16#07#),
      3849 => to_slv(opcode_type, 16#09#),
      3850 => to_slv(opcode_type, 16#0B#),
      3851 => to_slv(opcode_type, 16#0E#),
      3852 => to_slv(opcode_type, 16#06#),
      3853 => to_slv(opcode_type, 16#0F#),
      3854 => to_slv(opcode_type, 16#0F#),
      3855 => to_slv(opcode_type, 16#09#),
      3856 => to_slv(opcode_type, 16#06#),
      3857 => to_slv(opcode_type, 16#04#),
      3858 => to_slv(opcode_type, 16#21#),
      3859 => to_slv(opcode_type, 16#09#),
      3860 => to_slv(opcode_type, 16#11#),
      3861 => to_slv(opcode_type, 16#0D#),
      3862 => to_slv(opcode_type, 16#06#),
      3863 => to_slv(opcode_type, 16#07#),
      3864 => to_slv(opcode_type, 16#0C#),
      3865 => to_slv(opcode_type, 16#10#),
      3866 => to_slv(opcode_type, 16#07#),
      3867 => to_slv(opcode_type, 16#0D#),
      3868 => to_slv(opcode_type, 16#0B#),
      3869 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#07#),
      3873 => to_slv(opcode_type, 16#06#),
      3874 => to_slv(opcode_type, 16#09#),
      3875 => to_slv(opcode_type, 16#09#),
      3876 => to_slv(opcode_type, 16#11#),
      3877 => to_slv(opcode_type, 16#0B#),
      3878 => to_slv(opcode_type, 16#04#),
      3879 => to_slv(opcode_type, 16#10#),
      3880 => to_slv(opcode_type, 16#08#),
      3881 => to_slv(opcode_type, 16#06#),
      3882 => to_slv(opcode_type, 16#11#),
      3883 => to_slv(opcode_type, 16#0E#),
      3884 => to_slv(opcode_type, 16#09#),
      3885 => to_slv(opcode_type, 16#0B#),
      3886 => to_slv(opcode_type, 16#10#),
      3887 => to_slv(opcode_type, 16#09#),
      3888 => to_slv(opcode_type, 16#06#),
      3889 => to_slv(opcode_type, 16#03#),
      3890 => to_slv(opcode_type, 16#0C#),
      3891 => to_slv(opcode_type, 16#09#),
      3892 => to_slv(opcode_type, 16#0C#),
      3893 => to_slv(opcode_type, 16#11#),
      3894 => to_slv(opcode_type, 16#09#),
      3895 => to_slv(opcode_type, 16#08#),
      3896 => to_slv(opcode_type, 16#10#),
      3897 => to_slv(opcode_type, 16#10#),
      3898 => to_slv(opcode_type, 16#07#),
      3899 => to_slv(opcode_type, 16#0C#),
      3900 => to_slv(opcode_type, 16#0A#),
      3901 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#09#),
      3905 => to_slv(opcode_type, 16#08#),
      3906 => to_slv(opcode_type, 16#07#),
      3907 => to_slv(opcode_type, 16#09#),
      3908 => to_slv(opcode_type, 16#0D#),
      3909 => to_slv(opcode_type, 16#0A#),
      3910 => to_slv(opcode_type, 16#05#),
      3911 => to_slv(opcode_type, 16#10#),
      3912 => to_slv(opcode_type, 16#06#),
      3913 => to_slv(opcode_type, 16#05#),
      3914 => to_slv(opcode_type, 16#0B#),
      3915 => to_slv(opcode_type, 16#08#),
      3916 => to_slv(opcode_type, 16#0A#),
      3917 => to_slv(opcode_type, 16#0C#),
      3918 => to_slv(opcode_type, 16#08#),
      3919 => to_slv(opcode_type, 16#08#),
      3920 => to_slv(opcode_type, 16#08#),
      3921 => to_slv(opcode_type, 16#0A#),
      3922 => to_slv(opcode_type, 16#0A#),
      3923 => to_slv(opcode_type, 16#08#),
      3924 => to_slv(opcode_type, 16#0D#),
      3925 => to_slv(opcode_type, 16#0B#),
      3926 => to_slv(opcode_type, 16#08#),
      3927 => to_slv(opcode_type, 16#07#),
      3928 => to_slv(opcode_type, 16#0C#),
      3929 => to_slv(opcode_type, 16#0C#),
      3930 => to_slv(opcode_type, 16#07#),
      3931 => to_slv(opcode_type, 16#48#),
      3932 => to_slv(opcode_type, 16#31#),
      3933 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#09#),
      3937 => to_slv(opcode_type, 16#08#),
      3938 => to_slv(opcode_type, 16#07#),
      3939 => to_slv(opcode_type, 16#02#),
      3940 => to_slv(opcode_type, 16#0F#),
      3941 => to_slv(opcode_type, 16#07#),
      3942 => to_slv(opcode_type, 16#0F#),
      3943 => to_slv(opcode_type, 16#0D#),
      3944 => to_slv(opcode_type, 16#09#),
      3945 => to_slv(opcode_type, 16#01#),
      3946 => to_slv(opcode_type, 16#91#),
      3947 => to_slv(opcode_type, 16#06#),
      3948 => to_slv(opcode_type, 16#48#),
      3949 => to_slv(opcode_type, 16#0E#),
      3950 => to_slv(opcode_type, 16#06#),
      3951 => to_slv(opcode_type, 16#07#),
      3952 => to_slv(opcode_type, 16#08#),
      3953 => to_slv(opcode_type, 16#0B#),
      3954 => to_slv(opcode_type, 16#0C#),
      3955 => to_slv(opcode_type, 16#08#),
      3956 => to_slv(opcode_type, 16#74#),
      3957 => to_slv(opcode_type, 16#40#),
      3958 => to_slv(opcode_type, 16#09#),
      3959 => to_slv(opcode_type, 16#09#),
      3960 => to_slv(opcode_type, 16#0F#),
      3961 => to_slv(opcode_type, 16#0A#),
      3962 => to_slv(opcode_type, 16#08#),
      3963 => to_slv(opcode_type, 16#0A#),
      3964 => to_slv(opcode_type, 16#11#),
      3965 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#08#),
      3969 => to_slv(opcode_type, 16#09#),
      3970 => to_slv(opcode_type, 16#08#),
      3971 => to_slv(opcode_type, 16#07#),
      3972 => to_slv(opcode_type, 16#0D#),
      3973 => to_slv(opcode_type, 16#0B#),
      3974 => to_slv(opcode_type, 16#05#),
      3975 => to_slv(opcode_type, 16#11#),
      3976 => to_slv(opcode_type, 16#09#),
      3977 => to_slv(opcode_type, 16#06#),
      3978 => to_slv(opcode_type, 16#11#),
      3979 => to_slv(opcode_type, 16#0E#),
      3980 => to_slv(opcode_type, 16#02#),
      3981 => to_slv(opcode_type, 16#0D#),
      3982 => to_slv(opcode_type, 16#08#),
      3983 => to_slv(opcode_type, 16#06#),
      3984 => to_slv(opcode_type, 16#07#),
      3985 => to_slv(opcode_type, 16#0E#),
      3986 => to_slv(opcode_type, 16#11#),
      3987 => to_slv(opcode_type, 16#08#),
      3988 => to_slv(opcode_type, 16#11#),
      3989 => to_slv(opcode_type, 16#10#),
      3990 => to_slv(opcode_type, 16#08#),
      3991 => to_slv(opcode_type, 16#08#),
      3992 => to_slv(opcode_type, 16#0E#),
      3993 => to_slv(opcode_type, 16#0A#),
      3994 => to_slv(opcode_type, 16#07#),
      3995 => to_slv(opcode_type, 16#0C#),
      3996 => to_slv(opcode_type, 16#11#),
      3997 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#09#),
      4001 => to_slv(opcode_type, 16#08#),
      4002 => to_slv(opcode_type, 16#09#),
      4003 => to_slv(opcode_type, 16#03#),
      4004 => to_slv(opcode_type, 16#0A#),
      4005 => to_slv(opcode_type, 16#03#),
      4006 => to_slv(opcode_type, 16#10#),
      4007 => to_slv(opcode_type, 16#07#),
      4008 => to_slv(opcode_type, 16#06#),
      4009 => to_slv(opcode_type, 16#0D#),
      4010 => to_slv(opcode_type, 16#0C#),
      4011 => to_slv(opcode_type, 16#07#),
      4012 => to_slv(opcode_type, 16#0B#),
      4013 => to_slv(opcode_type, 16#0B#),
      4014 => to_slv(opcode_type, 16#09#),
      4015 => to_slv(opcode_type, 16#09#),
      4016 => to_slv(opcode_type, 16#09#),
      4017 => to_slv(opcode_type, 16#0A#),
      4018 => to_slv(opcode_type, 16#0B#),
      4019 => to_slv(opcode_type, 16#06#),
      4020 => to_slv(opcode_type, 16#0A#),
      4021 => to_slv(opcode_type, 16#0A#),
      4022 => to_slv(opcode_type, 16#06#),
      4023 => to_slv(opcode_type, 16#09#),
      4024 => to_slv(opcode_type, 16#0F#),
      4025 => to_slv(opcode_type, 16#0A#),
      4026 => to_slv(opcode_type, 16#06#),
      4027 => to_slv(opcode_type, 16#0D#),
      4028 => to_slv(opcode_type, 16#0B#),
      4029 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#06#),
      4033 => to_slv(opcode_type, 16#06#),
      4034 => to_slv(opcode_type, 16#06#),
      4035 => to_slv(opcode_type, 16#01#),
      4036 => to_slv(opcode_type, 16#11#),
      4037 => to_slv(opcode_type, 16#07#),
      4038 => to_slv(opcode_type, 16#79#),
      4039 => to_slv(opcode_type, 16#11#),
      4040 => to_slv(opcode_type, 16#06#),
      4041 => to_slv(opcode_type, 16#03#),
      4042 => to_slv(opcode_type, 16#0C#),
      4043 => to_slv(opcode_type, 16#07#),
      4044 => to_slv(opcode_type, 16#0D#),
      4045 => to_slv(opcode_type, 16#0B#),
      4046 => to_slv(opcode_type, 16#09#),
      4047 => to_slv(opcode_type, 16#09#),
      4048 => to_slv(opcode_type, 16#09#),
      4049 => to_slv(opcode_type, 16#0E#),
      4050 => to_slv(opcode_type, 16#E1#),
      4051 => to_slv(opcode_type, 16#09#),
      4052 => to_slv(opcode_type, 16#0D#),
      4053 => to_slv(opcode_type, 16#11#),
      4054 => to_slv(opcode_type, 16#09#),
      4055 => to_slv(opcode_type, 16#07#),
      4056 => to_slv(opcode_type, 16#10#),
      4057 => to_slv(opcode_type, 16#73#),
      4058 => to_slv(opcode_type, 16#07#),
      4059 => to_slv(opcode_type, 16#0F#),
      4060 => to_slv(opcode_type, 16#0B#),
      4061 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#08#),
      4065 => to_slv(opcode_type, 16#06#),
      4066 => to_slv(opcode_type, 16#09#),
      4067 => to_slv(opcode_type, 16#05#),
      4068 => to_slv(opcode_type, 16#0F#),
      4069 => to_slv(opcode_type, 16#07#),
      4070 => to_slv(opcode_type, 16#11#),
      4071 => to_slv(opcode_type, 16#11#),
      4072 => to_slv(opcode_type, 16#07#),
      4073 => to_slv(opcode_type, 16#06#),
      4074 => to_slv(opcode_type, 16#10#),
      4075 => to_slv(opcode_type, 16#0D#),
      4076 => to_slv(opcode_type, 16#06#),
      4077 => to_slv(opcode_type, 16#0E#),
      4078 => to_slv(opcode_type, 16#0B#),
      4079 => to_slv(opcode_type, 16#09#),
      4080 => to_slv(opcode_type, 16#09#),
      4081 => to_slv(opcode_type, 16#09#),
      4082 => to_slv(opcode_type, 16#0F#),
      4083 => to_slv(opcode_type, 16#0B#),
      4084 => to_slv(opcode_type, 16#07#),
      4085 => to_slv(opcode_type, 16#45#),
      4086 => to_slv(opcode_type, 16#0F#),
      4087 => to_slv(opcode_type, 16#07#),
      4088 => to_slv(opcode_type, 16#03#),
      4089 => to_slv(opcode_type, 16#0D#),
      4090 => to_slv(opcode_type, 16#09#),
      4091 => to_slv(opcode_type, 16#C7#),
      4092 => to_slv(opcode_type, 16#11#),
      4093 to 4095 => (others => '0')
  ),

    -- Bin `30`...
    29 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#06#),
      1 => to_slv(opcode_type, 16#06#),
      2 => to_slv(opcode_type, 16#08#),
      3 => to_slv(opcode_type, 16#01#),
      4 => to_slv(opcode_type, 16#0C#),
      5 => to_slv(opcode_type, 16#09#),
      6 => to_slv(opcode_type, 16#0A#),
      7 => to_slv(opcode_type, 16#10#),
      8 => to_slv(opcode_type, 16#08#),
      9 => to_slv(opcode_type, 16#07#),
      10 => to_slv(opcode_type, 16#0E#),
      11 => to_slv(opcode_type, 16#0F#),
      12 => to_slv(opcode_type, 16#08#),
      13 => to_slv(opcode_type, 16#72#),
      14 => to_slv(opcode_type, 16#0D#),
      15 => to_slv(opcode_type, 16#06#),
      16 => to_slv(opcode_type, 16#08#),
      17 => to_slv(opcode_type, 16#06#),
      18 => to_slv(opcode_type, 16#0E#),
      19 => to_slv(opcode_type, 16#0B#),
      20 => to_slv(opcode_type, 16#08#),
      21 => to_slv(opcode_type, 16#11#),
      22 => to_slv(opcode_type, 16#10#),
      23 => to_slv(opcode_type, 16#09#),
      24 => to_slv(opcode_type, 16#06#),
      25 => to_slv(opcode_type, 16#0B#),
      26 => to_slv(opcode_type, 16#7A#),
      27 => to_slv(opcode_type, 16#07#),
      28 => to_slv(opcode_type, 16#0E#),
      29 => to_slv(opcode_type, 16#59#),
      30 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#09#),
      33 => to_slv(opcode_type, 16#07#),
      34 => to_slv(opcode_type, 16#08#),
      35 => to_slv(opcode_type, 16#08#),
      36 => to_slv(opcode_type, 16#0B#),
      37 => to_slv(opcode_type, 16#0F#),
      38 => to_slv(opcode_type, 16#02#),
      39 => to_slv(opcode_type, 16#0A#),
      40 => to_slv(opcode_type, 16#07#),
      41 => to_slv(opcode_type, 16#08#),
      42 => to_slv(opcode_type, 16#0D#),
      43 => to_slv(opcode_type, 16#11#),
      44 => to_slv(opcode_type, 16#08#),
      45 => to_slv(opcode_type, 16#0B#),
      46 => to_slv(opcode_type, 16#0E#),
      47 => to_slv(opcode_type, 16#07#),
      48 => to_slv(opcode_type, 16#08#),
      49 => to_slv(opcode_type, 16#09#),
      50 => to_slv(opcode_type, 16#0E#),
      51 => to_slv(opcode_type, 16#11#),
      52 => to_slv(opcode_type, 16#07#),
      53 => to_slv(opcode_type, 16#0C#),
      54 => to_slv(opcode_type, 16#0D#),
      55 => to_slv(opcode_type, 16#09#),
      56 => to_slv(opcode_type, 16#07#),
      57 => to_slv(opcode_type, 16#10#),
      58 => to_slv(opcode_type, 16#10#),
      59 => to_slv(opcode_type, 16#09#),
      60 => to_slv(opcode_type, 16#10#),
      61 => to_slv(opcode_type, 16#0F#),
      62 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#09#),
      65 => to_slv(opcode_type, 16#07#),
      66 => to_slv(opcode_type, 16#09#),
      67 => to_slv(opcode_type, 16#05#),
      68 => to_slv(opcode_type, 16#1E#),
      69 => to_slv(opcode_type, 16#07#),
      70 => to_slv(opcode_type, 16#0D#),
      71 => to_slv(opcode_type, 16#0F#),
      72 => to_slv(opcode_type, 16#09#),
      73 => to_slv(opcode_type, 16#07#),
      74 => to_slv(opcode_type, 16#A6#),
      75 => to_slv(opcode_type, 16#0D#),
      76 => to_slv(opcode_type, 16#06#),
      77 => to_slv(opcode_type, 16#4E#),
      78 => to_slv(opcode_type, 16#10#),
      79 => to_slv(opcode_type, 16#08#),
      80 => to_slv(opcode_type, 16#06#),
      81 => to_slv(opcode_type, 16#09#),
      82 => to_slv(opcode_type, 16#97#),
      83 => to_slv(opcode_type, 16#11#),
      84 => to_slv(opcode_type, 16#06#),
      85 => to_slv(opcode_type, 16#11#),
      86 => to_slv(opcode_type, 16#11#),
      87 => to_slv(opcode_type, 16#07#),
      88 => to_slv(opcode_type, 16#06#),
      89 => to_slv(opcode_type, 16#0E#),
      90 => to_slv(opcode_type, 16#0C#),
      91 => to_slv(opcode_type, 16#09#),
      92 => to_slv(opcode_type, 16#11#),
      93 => to_slv(opcode_type, 16#A3#),
      94 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#06#),
      97 => to_slv(opcode_type, 16#09#),
      98 => to_slv(opcode_type, 16#08#),
      99 => to_slv(opcode_type, 16#08#),
      100 => to_slv(opcode_type, 16#0F#),
      101 => to_slv(opcode_type, 16#0E#),
      102 => to_slv(opcode_type, 16#06#),
      103 => to_slv(opcode_type, 16#0F#),
      104 => to_slv(opcode_type, 16#0C#),
      105 => to_slv(opcode_type, 16#07#),
      106 => to_slv(opcode_type, 16#07#),
      107 => to_slv(opcode_type, 16#0D#),
      108 => to_slv(opcode_type, 16#11#),
      109 => to_slv(opcode_type, 16#04#),
      110 => to_slv(opcode_type, 16#0E#),
      111 => to_slv(opcode_type, 16#07#),
      112 => to_slv(opcode_type, 16#09#),
      113 => to_slv(opcode_type, 16#09#),
      114 => to_slv(opcode_type, 16#31#),
      115 => to_slv(opcode_type, 16#0C#),
      116 => to_slv(opcode_type, 16#08#),
      117 => to_slv(opcode_type, 16#EA#),
      118 => to_slv(opcode_type, 16#11#),
      119 => to_slv(opcode_type, 16#06#),
      120 => to_slv(opcode_type, 16#09#),
      121 => to_slv(opcode_type, 16#0F#),
      122 => to_slv(opcode_type, 16#10#),
      123 => to_slv(opcode_type, 16#07#),
      124 => to_slv(opcode_type, 16#0A#),
      125 => to_slv(opcode_type, 16#0F#),
      126 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#07#),
      129 => to_slv(opcode_type, 16#06#),
      130 => to_slv(opcode_type, 16#06#),
      131 => to_slv(opcode_type, 16#03#),
      132 => to_slv(opcode_type, 16#0A#),
      133 => to_slv(opcode_type, 16#06#),
      134 => to_slv(opcode_type, 16#0D#),
      135 => to_slv(opcode_type, 16#0B#),
      136 => to_slv(opcode_type, 16#09#),
      137 => to_slv(opcode_type, 16#07#),
      138 => to_slv(opcode_type, 16#0A#),
      139 => to_slv(opcode_type, 16#0C#),
      140 => to_slv(opcode_type, 16#07#),
      141 => to_slv(opcode_type, 16#0F#),
      142 => to_slv(opcode_type, 16#11#),
      143 => to_slv(opcode_type, 16#06#),
      144 => to_slv(opcode_type, 16#07#),
      145 => to_slv(opcode_type, 16#08#),
      146 => to_slv(opcode_type, 16#10#),
      147 => to_slv(opcode_type, 16#0C#),
      148 => to_slv(opcode_type, 16#08#),
      149 => to_slv(opcode_type, 16#10#),
      150 => to_slv(opcode_type, 16#0A#),
      151 => to_slv(opcode_type, 16#08#),
      152 => to_slv(opcode_type, 16#06#),
      153 => to_slv(opcode_type, 16#0D#),
      154 => to_slv(opcode_type, 16#0D#),
      155 => to_slv(opcode_type, 16#06#),
      156 => to_slv(opcode_type, 16#0A#),
      157 => to_slv(opcode_type, 16#0C#),
      158 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#08#),
      161 => to_slv(opcode_type, 16#08#),
      162 => to_slv(opcode_type, 16#09#),
      163 => to_slv(opcode_type, 16#03#),
      164 => to_slv(opcode_type, 16#18#),
      165 => to_slv(opcode_type, 16#07#),
      166 => to_slv(opcode_type, 16#0E#),
      167 => to_slv(opcode_type, 16#13#),
      168 => to_slv(opcode_type, 16#07#),
      169 => to_slv(opcode_type, 16#08#),
      170 => to_slv(opcode_type, 16#11#),
      171 => to_slv(opcode_type, 16#0E#),
      172 => to_slv(opcode_type, 16#08#),
      173 => to_slv(opcode_type, 16#0D#),
      174 => to_slv(opcode_type, 16#0A#),
      175 => to_slv(opcode_type, 16#08#),
      176 => to_slv(opcode_type, 16#09#),
      177 => to_slv(opcode_type, 16#09#),
      178 => to_slv(opcode_type, 16#0A#),
      179 => to_slv(opcode_type, 16#86#),
      180 => to_slv(opcode_type, 16#09#),
      181 => to_slv(opcode_type, 16#0C#),
      182 => to_slv(opcode_type, 16#0A#),
      183 => to_slv(opcode_type, 16#06#),
      184 => to_slv(opcode_type, 16#06#),
      185 => to_slv(opcode_type, 16#0C#),
      186 => to_slv(opcode_type, 16#0F#),
      187 => to_slv(opcode_type, 16#08#),
      188 => to_slv(opcode_type, 16#0A#),
      189 => to_slv(opcode_type, 16#0E#),
      190 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#06#),
      193 => to_slv(opcode_type, 16#08#),
      194 => to_slv(opcode_type, 16#08#),
      195 => to_slv(opcode_type, 16#05#),
      196 => to_slv(opcode_type, 16#0E#),
      197 => to_slv(opcode_type, 16#08#),
      198 => to_slv(opcode_type, 16#0E#),
      199 => to_slv(opcode_type, 16#0D#),
      200 => to_slv(opcode_type, 16#07#),
      201 => to_slv(opcode_type, 16#08#),
      202 => to_slv(opcode_type, 16#0F#),
      203 => to_slv(opcode_type, 16#0A#),
      204 => to_slv(opcode_type, 16#06#),
      205 => to_slv(opcode_type, 16#0E#),
      206 => to_slv(opcode_type, 16#0C#),
      207 => to_slv(opcode_type, 16#09#),
      208 => to_slv(opcode_type, 16#08#),
      209 => to_slv(opcode_type, 16#07#),
      210 => to_slv(opcode_type, 16#10#),
      211 => to_slv(opcode_type, 16#0B#),
      212 => to_slv(opcode_type, 16#06#),
      213 => to_slv(opcode_type, 16#10#),
      214 => to_slv(opcode_type, 16#10#),
      215 => to_slv(opcode_type, 16#08#),
      216 => to_slv(opcode_type, 16#06#),
      217 => to_slv(opcode_type, 16#10#),
      218 => to_slv(opcode_type, 16#10#),
      219 => to_slv(opcode_type, 16#07#),
      220 => to_slv(opcode_type, 16#0E#),
      221 => to_slv(opcode_type, 16#0C#),
      222 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#07#),
      225 => to_slv(opcode_type, 16#08#),
      226 => to_slv(opcode_type, 16#07#),
      227 => to_slv(opcode_type, 16#07#),
      228 => to_slv(opcode_type, 16#10#),
      229 => to_slv(opcode_type, 16#0D#),
      230 => to_slv(opcode_type, 16#02#),
      231 => to_slv(opcode_type, 16#0A#),
      232 => to_slv(opcode_type, 16#07#),
      233 => to_slv(opcode_type, 16#07#),
      234 => to_slv(opcode_type, 16#0A#),
      235 => to_slv(opcode_type, 16#11#),
      236 => to_slv(opcode_type, 16#06#),
      237 => to_slv(opcode_type, 16#73#),
      238 => to_slv(opcode_type, 16#0E#),
      239 => to_slv(opcode_type, 16#06#),
      240 => to_slv(opcode_type, 16#07#),
      241 => to_slv(opcode_type, 16#07#),
      242 => to_slv(opcode_type, 16#0D#),
      243 => to_slv(opcode_type, 16#10#),
      244 => to_slv(opcode_type, 16#07#),
      245 => to_slv(opcode_type, 16#0E#),
      246 => to_slv(opcode_type, 16#0A#),
      247 => to_slv(opcode_type, 16#07#),
      248 => to_slv(opcode_type, 16#06#),
      249 => to_slv(opcode_type, 16#10#),
      250 => to_slv(opcode_type, 16#0D#),
      251 => to_slv(opcode_type, 16#08#),
      252 => to_slv(opcode_type, 16#82#),
      253 => to_slv(opcode_type, 16#0B#),
      254 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#06#),
      257 => to_slv(opcode_type, 16#07#),
      258 => to_slv(opcode_type, 16#09#),
      259 => to_slv(opcode_type, 16#07#),
      260 => to_slv(opcode_type, 16#10#),
      261 => to_slv(opcode_type, 16#10#),
      262 => to_slv(opcode_type, 16#06#),
      263 => to_slv(opcode_type, 16#0C#),
      264 => to_slv(opcode_type, 16#0F#),
      265 => to_slv(opcode_type, 16#07#),
      266 => to_slv(opcode_type, 16#08#),
      267 => to_slv(opcode_type, 16#0B#),
      268 => to_slv(opcode_type, 16#0F#),
      269 => to_slv(opcode_type, 16#01#),
      270 => to_slv(opcode_type, 16#0B#),
      271 => to_slv(opcode_type, 16#06#),
      272 => to_slv(opcode_type, 16#07#),
      273 => to_slv(opcode_type, 16#06#),
      274 => to_slv(opcode_type, 16#11#),
      275 => to_slv(opcode_type, 16#0A#),
      276 => to_slv(opcode_type, 16#09#),
      277 => to_slv(opcode_type, 16#11#),
      278 => to_slv(opcode_type, 16#0D#),
      279 => to_slv(opcode_type, 16#07#),
      280 => to_slv(opcode_type, 16#06#),
      281 => to_slv(opcode_type, 16#0A#),
      282 => to_slv(opcode_type, 16#0B#),
      283 => to_slv(opcode_type, 16#09#),
      284 => to_slv(opcode_type, 16#0C#),
      285 => to_slv(opcode_type, 16#0F#),
      286 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#09#),
      290 => to_slv(opcode_type, 16#08#),
      291 => to_slv(opcode_type, 16#09#),
      292 => to_slv(opcode_type, 16#0E#),
      293 => to_slv(opcode_type, 16#0E#),
      294 => to_slv(opcode_type, 16#07#),
      295 => to_slv(opcode_type, 16#FF#),
      296 => to_slv(opcode_type, 16#11#),
      297 => to_slv(opcode_type, 16#09#),
      298 => to_slv(opcode_type, 16#04#),
      299 => to_slv(opcode_type, 16#11#),
      300 => to_slv(opcode_type, 16#07#),
      301 => to_slv(opcode_type, 16#DB#),
      302 => to_slv(opcode_type, 16#0D#),
      303 => to_slv(opcode_type, 16#07#),
      304 => to_slv(opcode_type, 16#06#),
      305 => to_slv(opcode_type, 16#06#),
      306 => to_slv(opcode_type, 16#0E#),
      307 => to_slv(opcode_type, 16#0C#),
      308 => to_slv(opcode_type, 16#07#),
      309 => to_slv(opcode_type, 16#0A#),
      310 => to_slv(opcode_type, 16#11#),
      311 => to_slv(opcode_type, 16#08#),
      312 => to_slv(opcode_type, 16#06#),
      313 => to_slv(opcode_type, 16#0D#),
      314 => to_slv(opcode_type, 16#10#),
      315 => to_slv(opcode_type, 16#06#),
      316 => to_slv(opcode_type, 16#0A#),
      317 => to_slv(opcode_type, 16#0B#),
      318 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#07#),
      321 => to_slv(opcode_type, 16#08#),
      322 => to_slv(opcode_type, 16#09#),
      323 => to_slv(opcode_type, 16#07#),
      324 => to_slv(opcode_type, 16#0F#),
      325 => to_slv(opcode_type, 16#10#),
      326 => to_slv(opcode_type, 16#08#),
      327 => to_slv(opcode_type, 16#0F#),
      328 => to_slv(opcode_type, 16#75#),
      329 => to_slv(opcode_type, 16#08#),
      330 => to_slv(opcode_type, 16#06#),
      331 => to_slv(opcode_type, 16#0A#),
      332 => to_slv(opcode_type, 16#0B#),
      333 => to_slv(opcode_type, 16#01#),
      334 => to_slv(opcode_type, 16#11#),
      335 => to_slv(opcode_type, 16#07#),
      336 => to_slv(opcode_type, 16#06#),
      337 => to_slv(opcode_type, 16#08#),
      338 => to_slv(opcode_type, 16#0A#),
      339 => to_slv(opcode_type, 16#0E#),
      340 => to_slv(opcode_type, 16#09#),
      341 => to_slv(opcode_type, 16#E9#),
      342 => to_slv(opcode_type, 16#0C#),
      343 => to_slv(opcode_type, 16#06#),
      344 => to_slv(opcode_type, 16#07#),
      345 => to_slv(opcode_type, 16#11#),
      346 => to_slv(opcode_type, 16#10#),
      347 => to_slv(opcode_type, 16#07#),
      348 => to_slv(opcode_type, 16#0F#),
      349 => to_slv(opcode_type, 16#0E#),
      350 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#09#),
      353 => to_slv(opcode_type, 16#07#),
      354 => to_slv(opcode_type, 16#07#),
      355 => to_slv(opcode_type, 16#01#),
      356 => to_slv(opcode_type, 16#10#),
      357 => to_slv(opcode_type, 16#06#),
      358 => to_slv(opcode_type, 16#0D#),
      359 => to_slv(opcode_type, 16#0B#),
      360 => to_slv(opcode_type, 16#07#),
      361 => to_slv(opcode_type, 16#08#),
      362 => to_slv(opcode_type, 16#0B#),
      363 => to_slv(opcode_type, 16#0A#),
      364 => to_slv(opcode_type, 16#06#),
      365 => to_slv(opcode_type, 16#0A#),
      366 => to_slv(opcode_type, 16#0A#),
      367 => to_slv(opcode_type, 16#08#),
      368 => to_slv(opcode_type, 16#06#),
      369 => to_slv(opcode_type, 16#06#),
      370 => to_slv(opcode_type, 16#0B#),
      371 => to_slv(opcode_type, 16#0C#),
      372 => to_slv(opcode_type, 16#06#),
      373 => to_slv(opcode_type, 16#BD#),
      374 => to_slv(opcode_type, 16#D1#),
      375 => to_slv(opcode_type, 16#06#),
      376 => to_slv(opcode_type, 16#07#),
      377 => to_slv(opcode_type, 16#0E#),
      378 => to_slv(opcode_type, 16#0E#),
      379 => to_slv(opcode_type, 16#06#),
      380 => to_slv(opcode_type, 16#0C#),
      381 => to_slv(opcode_type, 16#0E#),
      382 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#07#),
      385 => to_slv(opcode_type, 16#09#),
      386 => to_slv(opcode_type, 16#07#),
      387 => to_slv(opcode_type, 16#04#),
      388 => to_slv(opcode_type, 16#B1#),
      389 => to_slv(opcode_type, 16#06#),
      390 => to_slv(opcode_type, 16#10#),
      391 => to_slv(opcode_type, 16#10#),
      392 => to_slv(opcode_type, 16#06#),
      393 => to_slv(opcode_type, 16#06#),
      394 => to_slv(opcode_type, 16#10#),
      395 => to_slv(opcode_type, 16#0E#),
      396 => to_slv(opcode_type, 16#06#),
      397 => to_slv(opcode_type, 16#0C#),
      398 => to_slv(opcode_type, 16#0F#),
      399 => to_slv(opcode_type, 16#06#),
      400 => to_slv(opcode_type, 16#06#),
      401 => to_slv(opcode_type, 16#08#),
      402 => to_slv(opcode_type, 16#0E#),
      403 => to_slv(opcode_type, 16#11#),
      404 => to_slv(opcode_type, 16#07#),
      405 => to_slv(opcode_type, 16#10#),
      406 => to_slv(opcode_type, 16#0B#),
      407 => to_slv(opcode_type, 16#08#),
      408 => to_slv(opcode_type, 16#07#),
      409 => to_slv(opcode_type, 16#11#),
      410 => to_slv(opcode_type, 16#70#),
      411 => to_slv(opcode_type, 16#08#),
      412 => to_slv(opcode_type, 16#0B#),
      413 => to_slv(opcode_type, 16#0E#),
      414 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#09#),
      417 => to_slv(opcode_type, 16#06#),
      418 => to_slv(opcode_type, 16#08#),
      419 => to_slv(opcode_type, 16#07#),
      420 => to_slv(opcode_type, 16#0B#),
      421 => to_slv(opcode_type, 16#11#),
      422 => to_slv(opcode_type, 16#08#),
      423 => to_slv(opcode_type, 16#0B#),
      424 => to_slv(opcode_type, 16#0D#),
      425 => to_slv(opcode_type, 16#07#),
      426 => to_slv(opcode_type, 16#01#),
      427 => to_slv(opcode_type, 16#0C#),
      428 => to_slv(opcode_type, 16#09#),
      429 => to_slv(opcode_type, 16#0C#),
      430 => to_slv(opcode_type, 16#11#),
      431 => to_slv(opcode_type, 16#06#),
      432 => to_slv(opcode_type, 16#06#),
      433 => to_slv(opcode_type, 16#07#),
      434 => to_slv(opcode_type, 16#0E#),
      435 => to_slv(opcode_type, 16#11#),
      436 => to_slv(opcode_type, 16#06#),
      437 => to_slv(opcode_type, 16#0C#),
      438 => to_slv(opcode_type, 16#11#),
      439 => to_slv(opcode_type, 16#08#),
      440 => to_slv(opcode_type, 16#08#),
      441 => to_slv(opcode_type, 16#0E#),
      442 => to_slv(opcode_type, 16#0D#),
      443 => to_slv(opcode_type, 16#08#),
      444 => to_slv(opcode_type, 16#11#),
      445 => to_slv(opcode_type, 16#0F#),
      446 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#08#),
      449 => to_slv(opcode_type, 16#09#),
      450 => to_slv(opcode_type, 16#06#),
      451 => to_slv(opcode_type, 16#08#),
      452 => to_slv(opcode_type, 16#0B#),
      453 => to_slv(opcode_type, 16#0E#),
      454 => to_slv(opcode_type, 16#02#),
      455 => to_slv(opcode_type, 16#0C#),
      456 => to_slv(opcode_type, 16#09#),
      457 => to_slv(opcode_type, 16#06#),
      458 => to_slv(opcode_type, 16#0C#),
      459 => to_slv(opcode_type, 16#5D#),
      460 => to_slv(opcode_type, 16#06#),
      461 => to_slv(opcode_type, 16#0C#),
      462 => to_slv(opcode_type, 16#10#),
      463 => to_slv(opcode_type, 16#06#),
      464 => to_slv(opcode_type, 16#09#),
      465 => to_slv(opcode_type, 16#08#),
      466 => to_slv(opcode_type, 16#11#),
      467 => to_slv(opcode_type, 16#0A#),
      468 => to_slv(opcode_type, 16#09#),
      469 => to_slv(opcode_type, 16#0E#),
      470 => to_slv(opcode_type, 16#0D#),
      471 => to_slv(opcode_type, 16#07#),
      472 => to_slv(opcode_type, 16#09#),
      473 => to_slv(opcode_type, 16#11#),
      474 => to_slv(opcode_type, 16#11#),
      475 => to_slv(opcode_type, 16#09#),
      476 => to_slv(opcode_type, 16#0E#),
      477 => to_slv(opcode_type, 16#0E#),
      478 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#07#),
      481 => to_slv(opcode_type, 16#06#),
      482 => to_slv(opcode_type, 16#08#),
      483 => to_slv(opcode_type, 16#01#),
      484 => to_slv(opcode_type, 16#0C#),
      485 => to_slv(opcode_type, 16#08#),
      486 => to_slv(opcode_type, 16#11#),
      487 => to_slv(opcode_type, 16#0D#),
      488 => to_slv(opcode_type, 16#08#),
      489 => to_slv(opcode_type, 16#09#),
      490 => to_slv(opcode_type, 16#0E#),
      491 => to_slv(opcode_type, 16#0A#),
      492 => to_slv(opcode_type, 16#08#),
      493 => to_slv(opcode_type, 16#11#),
      494 => to_slv(opcode_type, 16#0B#),
      495 => to_slv(opcode_type, 16#09#),
      496 => to_slv(opcode_type, 16#08#),
      497 => to_slv(opcode_type, 16#09#),
      498 => to_slv(opcode_type, 16#58#),
      499 => to_slv(opcode_type, 16#10#),
      500 => to_slv(opcode_type, 16#07#),
      501 => to_slv(opcode_type, 16#11#),
      502 => to_slv(opcode_type, 16#10#),
      503 => to_slv(opcode_type, 16#07#),
      504 => to_slv(opcode_type, 16#09#),
      505 => to_slv(opcode_type, 16#0C#),
      506 => to_slv(opcode_type, 16#0B#),
      507 => to_slv(opcode_type, 16#07#),
      508 => to_slv(opcode_type, 16#11#),
      509 => to_slv(opcode_type, 16#0A#),
      510 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#06#),
      513 => to_slv(opcode_type, 16#08#),
      514 => to_slv(opcode_type, 16#08#),
      515 => to_slv(opcode_type, 16#02#),
      516 => to_slv(opcode_type, 16#30#),
      517 => to_slv(opcode_type, 16#06#),
      518 => to_slv(opcode_type, 16#0B#),
      519 => to_slv(opcode_type, 16#10#),
      520 => to_slv(opcode_type, 16#09#),
      521 => to_slv(opcode_type, 16#07#),
      522 => to_slv(opcode_type, 16#10#),
      523 => to_slv(opcode_type, 16#0C#),
      524 => to_slv(opcode_type, 16#07#),
      525 => to_slv(opcode_type, 16#0F#),
      526 => to_slv(opcode_type, 16#11#),
      527 => to_slv(opcode_type, 16#07#),
      528 => to_slv(opcode_type, 16#07#),
      529 => to_slv(opcode_type, 16#06#),
      530 => to_slv(opcode_type, 16#0B#),
      531 => to_slv(opcode_type, 16#BA#),
      532 => to_slv(opcode_type, 16#08#),
      533 => to_slv(opcode_type, 16#0A#),
      534 => to_slv(opcode_type, 16#0E#),
      535 => to_slv(opcode_type, 16#08#),
      536 => to_slv(opcode_type, 16#06#),
      537 => to_slv(opcode_type, 16#10#),
      538 => to_slv(opcode_type, 16#84#),
      539 => to_slv(opcode_type, 16#06#),
      540 => to_slv(opcode_type, 16#AD#),
      541 => to_slv(opcode_type, 16#0B#),
      542 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#08#),
      545 => to_slv(opcode_type, 16#08#),
      546 => to_slv(opcode_type, 16#07#),
      547 => to_slv(opcode_type, 16#09#),
      548 => to_slv(opcode_type, 16#11#),
      549 => to_slv(opcode_type, 16#10#),
      550 => to_slv(opcode_type, 16#06#),
      551 => to_slv(opcode_type, 16#0F#),
      552 => to_slv(opcode_type, 16#0A#),
      553 => to_slv(opcode_type, 16#07#),
      554 => to_slv(opcode_type, 16#08#),
      555 => to_slv(opcode_type, 16#11#),
      556 => to_slv(opcode_type, 16#31#),
      557 => to_slv(opcode_type, 16#05#),
      558 => to_slv(opcode_type, 16#0B#),
      559 => to_slv(opcode_type, 16#09#),
      560 => to_slv(opcode_type, 16#07#),
      561 => to_slv(opcode_type, 16#06#),
      562 => to_slv(opcode_type, 16#0F#),
      563 => to_slv(opcode_type, 16#AA#),
      564 => to_slv(opcode_type, 16#09#),
      565 => to_slv(opcode_type, 16#0E#),
      566 => to_slv(opcode_type, 16#0C#),
      567 => to_slv(opcode_type, 16#07#),
      568 => to_slv(opcode_type, 16#07#),
      569 => to_slv(opcode_type, 16#11#),
      570 => to_slv(opcode_type, 16#0C#),
      571 => to_slv(opcode_type, 16#08#),
      572 => to_slv(opcode_type, 16#0E#),
      573 => to_slv(opcode_type, 16#0D#),
      574 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#06#),
      577 => to_slv(opcode_type, 16#06#),
      578 => to_slv(opcode_type, 16#07#),
      579 => to_slv(opcode_type, 16#07#),
      580 => to_slv(opcode_type, 16#0B#),
      581 => to_slv(opcode_type, 16#0B#),
      582 => to_slv(opcode_type, 16#06#),
      583 => to_slv(opcode_type, 16#0D#),
      584 => to_slv(opcode_type, 16#0A#),
      585 => to_slv(opcode_type, 16#09#),
      586 => to_slv(opcode_type, 16#06#),
      587 => to_slv(opcode_type, 16#10#),
      588 => to_slv(opcode_type, 16#0A#),
      589 => to_slv(opcode_type, 16#04#),
      590 => to_slv(opcode_type, 16#51#),
      591 => to_slv(opcode_type, 16#08#),
      592 => to_slv(opcode_type, 16#09#),
      593 => to_slv(opcode_type, 16#09#),
      594 => to_slv(opcode_type, 16#0C#),
      595 => to_slv(opcode_type, 16#0A#),
      596 => to_slv(opcode_type, 16#09#),
      597 => to_slv(opcode_type, 16#0A#),
      598 => to_slv(opcode_type, 16#10#),
      599 => to_slv(opcode_type, 16#08#),
      600 => to_slv(opcode_type, 16#09#),
      601 => to_slv(opcode_type, 16#0C#),
      602 => to_slv(opcode_type, 16#0D#),
      603 => to_slv(opcode_type, 16#09#),
      604 => to_slv(opcode_type, 16#11#),
      605 => to_slv(opcode_type, 16#11#),
      606 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#06#),
      609 => to_slv(opcode_type, 16#09#),
      610 => to_slv(opcode_type, 16#08#),
      611 => to_slv(opcode_type, 16#05#),
      612 => to_slv(opcode_type, 16#0E#),
      613 => to_slv(opcode_type, 16#07#),
      614 => to_slv(opcode_type, 16#10#),
      615 => to_slv(opcode_type, 16#0B#),
      616 => to_slv(opcode_type, 16#07#),
      617 => to_slv(opcode_type, 16#07#),
      618 => to_slv(opcode_type, 16#0E#),
      619 => to_slv(opcode_type, 16#68#),
      620 => to_slv(opcode_type, 16#07#),
      621 => to_slv(opcode_type, 16#0F#),
      622 => to_slv(opcode_type, 16#0E#),
      623 => to_slv(opcode_type, 16#09#),
      624 => to_slv(opcode_type, 16#07#),
      625 => to_slv(opcode_type, 16#08#),
      626 => to_slv(opcode_type, 16#0F#),
      627 => to_slv(opcode_type, 16#0D#),
      628 => to_slv(opcode_type, 16#07#),
      629 => to_slv(opcode_type, 16#11#),
      630 => to_slv(opcode_type, 16#10#),
      631 => to_slv(opcode_type, 16#07#),
      632 => to_slv(opcode_type, 16#08#),
      633 => to_slv(opcode_type, 16#10#),
      634 => to_slv(opcode_type, 16#11#),
      635 => to_slv(opcode_type, 16#09#),
      636 => to_slv(opcode_type, 16#0C#),
      637 => to_slv(opcode_type, 16#0B#),
      638 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#08#),
      641 => to_slv(opcode_type, 16#08#),
      642 => to_slv(opcode_type, 16#06#),
      643 => to_slv(opcode_type, 16#08#),
      644 => to_slv(opcode_type, 16#0F#),
      645 => to_slv(opcode_type, 16#6E#),
      646 => to_slv(opcode_type, 16#02#),
      647 => to_slv(opcode_type, 16#0D#),
      648 => to_slv(opcode_type, 16#07#),
      649 => to_slv(opcode_type, 16#09#),
      650 => to_slv(opcode_type, 16#10#),
      651 => to_slv(opcode_type, 16#0C#),
      652 => to_slv(opcode_type, 16#07#),
      653 => to_slv(opcode_type, 16#0C#),
      654 => to_slv(opcode_type, 16#0B#),
      655 => to_slv(opcode_type, 16#08#),
      656 => to_slv(opcode_type, 16#07#),
      657 => to_slv(opcode_type, 16#08#),
      658 => to_slv(opcode_type, 16#10#),
      659 => to_slv(opcode_type, 16#0E#),
      660 => to_slv(opcode_type, 16#06#),
      661 => to_slv(opcode_type, 16#0B#),
      662 => to_slv(opcode_type, 16#0C#),
      663 => to_slv(opcode_type, 16#07#),
      664 => to_slv(opcode_type, 16#06#),
      665 => to_slv(opcode_type, 16#0B#),
      666 => to_slv(opcode_type, 16#10#),
      667 => to_slv(opcode_type, 16#08#),
      668 => to_slv(opcode_type, 16#0F#),
      669 => to_slv(opcode_type, 16#0A#),
      670 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#09#),
      673 => to_slv(opcode_type, 16#06#),
      674 => to_slv(opcode_type, 16#09#),
      675 => to_slv(opcode_type, 16#04#),
      676 => to_slv(opcode_type, 16#10#),
      677 => to_slv(opcode_type, 16#07#),
      678 => to_slv(opcode_type, 16#0E#),
      679 => to_slv(opcode_type, 16#0B#),
      680 => to_slv(opcode_type, 16#07#),
      681 => to_slv(opcode_type, 16#07#),
      682 => to_slv(opcode_type, 16#11#),
      683 => to_slv(opcode_type, 16#0E#),
      684 => to_slv(opcode_type, 16#09#),
      685 => to_slv(opcode_type, 16#0F#),
      686 => to_slv(opcode_type, 16#0F#),
      687 => to_slv(opcode_type, 16#08#),
      688 => to_slv(opcode_type, 16#08#),
      689 => to_slv(opcode_type, 16#09#),
      690 => to_slv(opcode_type, 16#0B#),
      691 => to_slv(opcode_type, 16#0C#),
      692 => to_slv(opcode_type, 16#06#),
      693 => to_slv(opcode_type, 16#0A#),
      694 => to_slv(opcode_type, 16#11#),
      695 => to_slv(opcode_type, 16#09#),
      696 => to_slv(opcode_type, 16#06#),
      697 => to_slv(opcode_type, 16#0A#),
      698 => to_slv(opcode_type, 16#11#),
      699 => to_slv(opcode_type, 16#08#),
      700 => to_slv(opcode_type, 16#0F#),
      701 => to_slv(opcode_type, 16#0E#),
      702 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#08#),
      705 => to_slv(opcode_type, 16#09#),
      706 => to_slv(opcode_type, 16#06#),
      707 => to_slv(opcode_type, 16#05#),
      708 => to_slv(opcode_type, 16#11#),
      709 => to_slv(opcode_type, 16#06#),
      710 => to_slv(opcode_type, 16#11#),
      711 => to_slv(opcode_type, 16#0F#),
      712 => to_slv(opcode_type, 16#06#),
      713 => to_slv(opcode_type, 16#08#),
      714 => to_slv(opcode_type, 16#0B#),
      715 => to_slv(opcode_type, 16#FC#),
      716 => to_slv(opcode_type, 16#06#),
      717 => to_slv(opcode_type, 16#11#),
      718 => to_slv(opcode_type, 16#0F#),
      719 => to_slv(opcode_type, 16#06#),
      720 => to_slv(opcode_type, 16#09#),
      721 => to_slv(opcode_type, 16#09#),
      722 => to_slv(opcode_type, 16#11#),
      723 => to_slv(opcode_type, 16#0E#),
      724 => to_slv(opcode_type, 16#06#),
      725 => to_slv(opcode_type, 16#0F#),
      726 => to_slv(opcode_type, 16#0D#),
      727 => to_slv(opcode_type, 16#08#),
      728 => to_slv(opcode_type, 16#09#),
      729 => to_slv(opcode_type, 16#A2#),
      730 => to_slv(opcode_type, 16#10#),
      731 => to_slv(opcode_type, 16#06#),
      732 => to_slv(opcode_type, 16#11#),
      733 => to_slv(opcode_type, 16#0C#),
      734 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#07#),
      737 => to_slv(opcode_type, 16#09#),
      738 => to_slv(opcode_type, 16#06#),
      739 => to_slv(opcode_type, 16#04#),
      740 => to_slv(opcode_type, 16#0D#),
      741 => to_slv(opcode_type, 16#06#),
      742 => to_slv(opcode_type, 16#0C#),
      743 => to_slv(opcode_type, 16#10#),
      744 => to_slv(opcode_type, 16#08#),
      745 => to_slv(opcode_type, 16#07#),
      746 => to_slv(opcode_type, 16#0E#),
      747 => to_slv(opcode_type, 16#0C#),
      748 => to_slv(opcode_type, 16#08#),
      749 => to_slv(opcode_type, 16#0D#),
      750 => to_slv(opcode_type, 16#10#),
      751 => to_slv(opcode_type, 16#09#),
      752 => to_slv(opcode_type, 16#07#),
      753 => to_slv(opcode_type, 16#07#),
      754 => to_slv(opcode_type, 16#0C#),
      755 => to_slv(opcode_type, 16#0E#),
      756 => to_slv(opcode_type, 16#07#),
      757 => to_slv(opcode_type, 16#0B#),
      758 => to_slv(opcode_type, 16#10#),
      759 => to_slv(opcode_type, 16#09#),
      760 => to_slv(opcode_type, 16#07#),
      761 => to_slv(opcode_type, 16#0F#),
      762 => to_slv(opcode_type, 16#0A#),
      763 => to_slv(opcode_type, 16#06#),
      764 => to_slv(opcode_type, 16#0C#),
      765 => to_slv(opcode_type, 16#0E#),
      766 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#06#),
      769 => to_slv(opcode_type, 16#07#),
      770 => to_slv(opcode_type, 16#06#),
      771 => to_slv(opcode_type, 16#04#),
      772 => to_slv(opcode_type, 16#0C#),
      773 => to_slv(opcode_type, 16#08#),
      774 => to_slv(opcode_type, 16#11#),
      775 => to_slv(opcode_type, 16#0E#),
      776 => to_slv(opcode_type, 16#06#),
      777 => to_slv(opcode_type, 16#07#),
      778 => to_slv(opcode_type, 16#0D#),
      779 => to_slv(opcode_type, 16#10#),
      780 => to_slv(opcode_type, 16#07#),
      781 => to_slv(opcode_type, 16#0A#),
      782 => to_slv(opcode_type, 16#4C#),
      783 => to_slv(opcode_type, 16#08#),
      784 => to_slv(opcode_type, 16#09#),
      785 => to_slv(opcode_type, 16#09#),
      786 => to_slv(opcode_type, 16#11#),
      787 => to_slv(opcode_type, 16#DE#),
      788 => to_slv(opcode_type, 16#08#),
      789 => to_slv(opcode_type, 16#10#),
      790 => to_slv(opcode_type, 16#0A#),
      791 => to_slv(opcode_type, 16#06#),
      792 => to_slv(opcode_type, 16#07#),
      793 => to_slv(opcode_type, 16#0A#),
      794 => to_slv(opcode_type, 16#0E#),
      795 => to_slv(opcode_type, 16#08#),
      796 => to_slv(opcode_type, 16#0D#),
      797 => to_slv(opcode_type, 16#0A#),
      798 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#07#),
      801 => to_slv(opcode_type, 16#09#),
      802 => to_slv(opcode_type, 16#09#),
      803 => to_slv(opcode_type, 16#04#),
      804 => to_slv(opcode_type, 16#0A#),
      805 => to_slv(opcode_type, 16#08#),
      806 => to_slv(opcode_type, 16#0C#),
      807 => to_slv(opcode_type, 16#11#),
      808 => to_slv(opcode_type, 16#08#),
      809 => to_slv(opcode_type, 16#08#),
      810 => to_slv(opcode_type, 16#6D#),
      811 => to_slv(opcode_type, 16#0A#),
      812 => to_slv(opcode_type, 16#09#),
      813 => to_slv(opcode_type, 16#0A#),
      814 => to_slv(opcode_type, 16#0E#),
      815 => to_slv(opcode_type, 16#07#),
      816 => to_slv(opcode_type, 16#06#),
      817 => to_slv(opcode_type, 16#08#),
      818 => to_slv(opcode_type, 16#0A#),
      819 => to_slv(opcode_type, 16#11#),
      820 => to_slv(opcode_type, 16#09#),
      821 => to_slv(opcode_type, 16#11#),
      822 => to_slv(opcode_type, 16#0A#),
      823 => to_slv(opcode_type, 16#06#),
      824 => to_slv(opcode_type, 16#07#),
      825 => to_slv(opcode_type, 16#0C#),
      826 => to_slv(opcode_type, 16#0F#),
      827 => to_slv(opcode_type, 16#06#),
      828 => to_slv(opcode_type, 16#0A#),
      829 => to_slv(opcode_type, 16#0E#),
      830 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#06#),
      833 => to_slv(opcode_type, 16#06#),
      834 => to_slv(opcode_type, 16#06#),
      835 => to_slv(opcode_type, 16#01#),
      836 => to_slv(opcode_type, 16#28#),
      837 => to_slv(opcode_type, 16#06#),
      838 => to_slv(opcode_type, 16#0D#),
      839 => to_slv(opcode_type, 16#0A#),
      840 => to_slv(opcode_type, 16#09#),
      841 => to_slv(opcode_type, 16#06#),
      842 => to_slv(opcode_type, 16#0E#),
      843 => to_slv(opcode_type, 16#0E#),
      844 => to_slv(opcode_type, 16#08#),
      845 => to_slv(opcode_type, 16#0C#),
      846 => to_slv(opcode_type, 16#0A#),
      847 => to_slv(opcode_type, 16#07#),
      848 => to_slv(opcode_type, 16#06#),
      849 => to_slv(opcode_type, 16#08#),
      850 => to_slv(opcode_type, 16#E1#),
      851 => to_slv(opcode_type, 16#11#),
      852 => to_slv(opcode_type, 16#08#),
      853 => to_slv(opcode_type, 16#0F#),
      854 => to_slv(opcode_type, 16#0D#),
      855 => to_slv(opcode_type, 16#06#),
      856 => to_slv(opcode_type, 16#08#),
      857 => to_slv(opcode_type, 16#11#),
      858 => to_slv(opcode_type, 16#0A#),
      859 => to_slv(opcode_type, 16#06#),
      860 => to_slv(opcode_type, 16#11#),
      861 => to_slv(opcode_type, 16#0F#),
      862 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#07#),
      865 => to_slv(opcode_type, 16#07#),
      866 => to_slv(opcode_type, 16#07#),
      867 => to_slv(opcode_type, 16#06#),
      868 => to_slv(opcode_type, 16#0A#),
      869 => to_slv(opcode_type, 16#E4#),
      870 => to_slv(opcode_type, 16#08#),
      871 => to_slv(opcode_type, 16#0D#),
      872 => to_slv(opcode_type, 16#0D#),
      873 => to_slv(opcode_type, 16#07#),
      874 => to_slv(opcode_type, 16#01#),
      875 => to_slv(opcode_type, 16#11#),
      876 => to_slv(opcode_type, 16#08#),
      877 => to_slv(opcode_type, 16#67#),
      878 => to_slv(opcode_type, 16#B7#),
      879 => to_slv(opcode_type, 16#06#),
      880 => to_slv(opcode_type, 16#08#),
      881 => to_slv(opcode_type, 16#06#),
      882 => to_slv(opcode_type, 16#C3#),
      883 => to_slv(opcode_type, 16#0E#),
      884 => to_slv(opcode_type, 16#07#),
      885 => to_slv(opcode_type, 16#0B#),
      886 => to_slv(opcode_type, 16#0A#),
      887 => to_slv(opcode_type, 16#06#),
      888 => to_slv(opcode_type, 16#07#),
      889 => to_slv(opcode_type, 16#11#),
      890 => to_slv(opcode_type, 16#0A#),
      891 => to_slv(opcode_type, 16#07#),
      892 => to_slv(opcode_type, 16#0E#),
      893 => to_slv(opcode_type, 16#0B#),
      894 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#06#),
      897 => to_slv(opcode_type, 16#07#),
      898 => to_slv(opcode_type, 16#08#),
      899 => to_slv(opcode_type, 16#06#),
      900 => to_slv(opcode_type, 16#35#),
      901 => to_slv(opcode_type, 16#0C#),
      902 => to_slv(opcode_type, 16#06#),
      903 => to_slv(opcode_type, 16#11#),
      904 => to_slv(opcode_type, 16#0F#),
      905 => to_slv(opcode_type, 16#09#),
      906 => to_slv(opcode_type, 16#03#),
      907 => to_slv(opcode_type, 16#0B#),
      908 => to_slv(opcode_type, 16#09#),
      909 => to_slv(opcode_type, 16#11#),
      910 => to_slv(opcode_type, 16#0B#),
      911 => to_slv(opcode_type, 16#08#),
      912 => to_slv(opcode_type, 16#08#),
      913 => to_slv(opcode_type, 16#08#),
      914 => to_slv(opcode_type, 16#10#),
      915 => to_slv(opcode_type, 16#11#),
      916 => to_slv(opcode_type, 16#06#),
      917 => to_slv(opcode_type, 16#0A#),
      918 => to_slv(opcode_type, 16#0D#),
      919 => to_slv(opcode_type, 16#09#),
      920 => to_slv(opcode_type, 16#09#),
      921 => to_slv(opcode_type, 16#0A#),
      922 => to_slv(opcode_type, 16#11#),
      923 => to_slv(opcode_type, 16#08#),
      924 => to_slv(opcode_type, 16#0B#),
      925 => to_slv(opcode_type, 16#0C#),
      926 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#07#),
      929 => to_slv(opcode_type, 16#06#),
      930 => to_slv(opcode_type, 16#09#),
      931 => to_slv(opcode_type, 16#01#),
      932 => to_slv(opcode_type, 16#10#),
      933 => to_slv(opcode_type, 16#09#),
      934 => to_slv(opcode_type, 16#0D#),
      935 => to_slv(opcode_type, 16#0F#),
      936 => to_slv(opcode_type, 16#07#),
      937 => to_slv(opcode_type, 16#07#),
      938 => to_slv(opcode_type, 16#0E#),
      939 => to_slv(opcode_type, 16#0C#),
      940 => to_slv(opcode_type, 16#06#),
      941 => to_slv(opcode_type, 16#0F#),
      942 => to_slv(opcode_type, 16#0A#),
      943 => to_slv(opcode_type, 16#09#),
      944 => to_slv(opcode_type, 16#06#),
      945 => to_slv(opcode_type, 16#07#),
      946 => to_slv(opcode_type, 16#11#),
      947 => to_slv(opcode_type, 16#0E#),
      948 => to_slv(opcode_type, 16#09#),
      949 => to_slv(opcode_type, 16#0E#),
      950 => to_slv(opcode_type, 16#0E#),
      951 => to_slv(opcode_type, 16#06#),
      952 => to_slv(opcode_type, 16#06#),
      953 => to_slv(opcode_type, 16#1E#),
      954 => to_slv(opcode_type, 16#0A#),
      955 => to_slv(opcode_type, 16#08#),
      956 => to_slv(opcode_type, 16#0A#),
      957 => to_slv(opcode_type, 16#11#),
      958 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#07#),
      961 => to_slv(opcode_type, 16#06#),
      962 => to_slv(opcode_type, 16#09#),
      963 => to_slv(opcode_type, 16#05#),
      964 => to_slv(opcode_type, 16#0A#),
      965 => to_slv(opcode_type, 16#07#),
      966 => to_slv(opcode_type, 16#10#),
      967 => to_slv(opcode_type, 16#0A#),
      968 => to_slv(opcode_type, 16#06#),
      969 => to_slv(opcode_type, 16#06#),
      970 => to_slv(opcode_type, 16#76#),
      971 => to_slv(opcode_type, 16#10#),
      972 => to_slv(opcode_type, 16#07#),
      973 => to_slv(opcode_type, 16#0B#),
      974 => to_slv(opcode_type, 16#0F#),
      975 => to_slv(opcode_type, 16#07#),
      976 => to_slv(opcode_type, 16#09#),
      977 => to_slv(opcode_type, 16#07#),
      978 => to_slv(opcode_type, 16#0D#),
      979 => to_slv(opcode_type, 16#0E#),
      980 => to_slv(opcode_type, 16#07#),
      981 => to_slv(opcode_type, 16#11#),
      982 => to_slv(opcode_type, 16#0F#),
      983 => to_slv(opcode_type, 16#07#),
      984 => to_slv(opcode_type, 16#09#),
      985 => to_slv(opcode_type, 16#0E#),
      986 => to_slv(opcode_type, 16#0F#),
      987 => to_slv(opcode_type, 16#06#),
      988 => to_slv(opcode_type, 16#0E#),
      989 => to_slv(opcode_type, 16#0B#),
      990 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#06#),
      993 => to_slv(opcode_type, 16#09#),
      994 => to_slv(opcode_type, 16#08#),
      995 => to_slv(opcode_type, 16#04#),
      996 => to_slv(opcode_type, 16#0D#),
      997 => to_slv(opcode_type, 16#06#),
      998 => to_slv(opcode_type, 16#0E#),
      999 => to_slv(opcode_type, 16#0C#),
      1000 => to_slv(opcode_type, 16#06#),
      1001 => to_slv(opcode_type, 16#08#),
      1002 => to_slv(opcode_type, 16#0B#),
      1003 => to_slv(opcode_type, 16#0B#),
      1004 => to_slv(opcode_type, 16#06#),
      1005 => to_slv(opcode_type, 16#0F#),
      1006 => to_slv(opcode_type, 16#11#),
      1007 => to_slv(opcode_type, 16#08#),
      1008 => to_slv(opcode_type, 16#07#),
      1009 => to_slv(opcode_type, 16#08#),
      1010 => to_slv(opcode_type, 16#11#),
      1011 => to_slv(opcode_type, 16#0E#),
      1012 => to_slv(opcode_type, 16#09#),
      1013 => to_slv(opcode_type, 16#0B#),
      1014 => to_slv(opcode_type, 16#0D#),
      1015 => to_slv(opcode_type, 16#08#),
      1016 => to_slv(opcode_type, 16#06#),
      1017 => to_slv(opcode_type, 16#0B#),
      1018 => to_slv(opcode_type, 16#0C#),
      1019 => to_slv(opcode_type, 16#07#),
      1020 => to_slv(opcode_type, 16#12#),
      1021 => to_slv(opcode_type, 16#0E#),
      1022 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#06#),
      1025 => to_slv(opcode_type, 16#06#),
      1026 => to_slv(opcode_type, 16#09#),
      1027 => to_slv(opcode_type, 16#04#),
      1028 => to_slv(opcode_type, 16#0D#),
      1029 => to_slv(opcode_type, 16#07#),
      1030 => to_slv(opcode_type, 16#0C#),
      1031 => to_slv(opcode_type, 16#0D#),
      1032 => to_slv(opcode_type, 16#06#),
      1033 => to_slv(opcode_type, 16#08#),
      1034 => to_slv(opcode_type, 16#0A#),
      1035 => to_slv(opcode_type, 16#0A#),
      1036 => to_slv(opcode_type, 16#07#),
      1037 => to_slv(opcode_type, 16#0C#),
      1038 => to_slv(opcode_type, 16#0A#),
      1039 => to_slv(opcode_type, 16#06#),
      1040 => to_slv(opcode_type, 16#06#),
      1041 => to_slv(opcode_type, 16#09#),
      1042 => to_slv(opcode_type, 16#0A#),
      1043 => to_slv(opcode_type, 16#0C#),
      1044 => to_slv(opcode_type, 16#06#),
      1045 => to_slv(opcode_type, 16#11#),
      1046 => to_slv(opcode_type, 16#0F#),
      1047 => to_slv(opcode_type, 16#09#),
      1048 => to_slv(opcode_type, 16#09#),
      1049 => to_slv(opcode_type, 16#0C#),
      1050 => to_slv(opcode_type, 16#0D#),
      1051 => to_slv(opcode_type, 16#07#),
      1052 => to_slv(opcode_type, 16#0B#),
      1053 => to_slv(opcode_type, 16#0C#),
      1054 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#07#),
      1057 => to_slv(opcode_type, 16#09#),
      1058 => to_slv(opcode_type, 16#07#),
      1059 => to_slv(opcode_type, 16#05#),
      1060 => to_slv(opcode_type, 16#11#),
      1061 => to_slv(opcode_type, 16#08#),
      1062 => to_slv(opcode_type, 16#11#),
      1063 => to_slv(opcode_type, 16#10#),
      1064 => to_slv(opcode_type, 16#08#),
      1065 => to_slv(opcode_type, 16#08#),
      1066 => to_slv(opcode_type, 16#0C#),
      1067 => to_slv(opcode_type, 16#10#),
      1068 => to_slv(opcode_type, 16#07#),
      1069 => to_slv(opcode_type, 16#11#),
      1070 => to_slv(opcode_type, 16#0B#),
      1071 => to_slv(opcode_type, 16#07#),
      1072 => to_slv(opcode_type, 16#06#),
      1073 => to_slv(opcode_type, 16#06#),
      1074 => to_slv(opcode_type, 16#0A#),
      1075 => to_slv(opcode_type, 16#0E#),
      1076 => to_slv(opcode_type, 16#07#),
      1077 => to_slv(opcode_type, 16#0D#),
      1078 => to_slv(opcode_type, 16#11#),
      1079 => to_slv(opcode_type, 16#07#),
      1080 => to_slv(opcode_type, 16#08#),
      1081 => to_slv(opcode_type, 16#50#),
      1082 => to_slv(opcode_type, 16#0B#),
      1083 => to_slv(opcode_type, 16#08#),
      1084 => to_slv(opcode_type, 16#11#),
      1085 => to_slv(opcode_type, 16#0F#),
      1086 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#06#),
      1089 => to_slv(opcode_type, 16#07#),
      1090 => to_slv(opcode_type, 16#08#),
      1091 => to_slv(opcode_type, 16#08#),
      1092 => to_slv(opcode_type, 16#0C#),
      1093 => to_slv(opcode_type, 16#85#),
      1094 => to_slv(opcode_type, 16#05#),
      1095 => to_slv(opcode_type, 16#8D#),
      1096 => to_slv(opcode_type, 16#09#),
      1097 => to_slv(opcode_type, 16#06#),
      1098 => to_slv(opcode_type, 16#11#),
      1099 => to_slv(opcode_type, 16#0F#),
      1100 => to_slv(opcode_type, 16#09#),
      1101 => to_slv(opcode_type, 16#0B#),
      1102 => to_slv(opcode_type, 16#0A#),
      1103 => to_slv(opcode_type, 16#07#),
      1104 => to_slv(opcode_type, 16#08#),
      1105 => to_slv(opcode_type, 16#07#),
      1106 => to_slv(opcode_type, 16#0D#),
      1107 => to_slv(opcode_type, 16#0C#),
      1108 => to_slv(opcode_type, 16#07#),
      1109 => to_slv(opcode_type, 16#0F#),
      1110 => to_slv(opcode_type, 16#0A#),
      1111 => to_slv(opcode_type, 16#07#),
      1112 => to_slv(opcode_type, 16#08#),
      1113 => to_slv(opcode_type, 16#11#),
      1114 => to_slv(opcode_type, 16#C4#),
      1115 => to_slv(opcode_type, 16#06#),
      1116 => to_slv(opcode_type, 16#10#),
      1117 => to_slv(opcode_type, 16#0C#),
      1118 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#06#),
      1121 => to_slv(opcode_type, 16#07#),
      1122 => to_slv(opcode_type, 16#07#),
      1123 => to_slv(opcode_type, 16#07#),
      1124 => to_slv(opcode_type, 16#0D#),
      1125 => to_slv(opcode_type, 16#0F#),
      1126 => to_slv(opcode_type, 16#06#),
      1127 => to_slv(opcode_type, 16#11#),
      1128 => to_slv(opcode_type, 16#11#),
      1129 => to_slv(opcode_type, 16#09#),
      1130 => to_slv(opcode_type, 16#03#),
      1131 => to_slv(opcode_type, 16#0C#),
      1132 => to_slv(opcode_type, 16#08#),
      1133 => to_slv(opcode_type, 16#11#),
      1134 => to_slv(opcode_type, 16#0E#),
      1135 => to_slv(opcode_type, 16#09#),
      1136 => to_slv(opcode_type, 16#08#),
      1137 => to_slv(opcode_type, 16#06#),
      1138 => to_slv(opcode_type, 16#0F#),
      1139 => to_slv(opcode_type, 16#10#),
      1140 => to_slv(opcode_type, 16#09#),
      1141 => to_slv(opcode_type, 16#0A#),
      1142 => to_slv(opcode_type, 16#11#),
      1143 => to_slv(opcode_type, 16#09#),
      1144 => to_slv(opcode_type, 16#09#),
      1145 => to_slv(opcode_type, 16#0D#),
      1146 => to_slv(opcode_type, 16#0F#),
      1147 => to_slv(opcode_type, 16#07#),
      1148 => to_slv(opcode_type, 16#0D#),
      1149 => to_slv(opcode_type, 16#0F#),
      1150 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#07#),
      1153 => to_slv(opcode_type, 16#09#),
      1154 => to_slv(opcode_type, 16#08#),
      1155 => to_slv(opcode_type, 16#08#),
      1156 => to_slv(opcode_type, 16#0C#),
      1157 => to_slv(opcode_type, 16#D7#),
      1158 => to_slv(opcode_type, 16#01#),
      1159 => to_slv(opcode_type, 16#7A#),
      1160 => to_slv(opcode_type, 16#09#),
      1161 => to_slv(opcode_type, 16#09#),
      1162 => to_slv(opcode_type, 16#0E#),
      1163 => to_slv(opcode_type, 16#65#),
      1164 => to_slv(opcode_type, 16#09#),
      1165 => to_slv(opcode_type, 16#11#),
      1166 => to_slv(opcode_type, 16#0F#),
      1167 => to_slv(opcode_type, 16#06#),
      1168 => to_slv(opcode_type, 16#06#),
      1169 => to_slv(opcode_type, 16#07#),
      1170 => to_slv(opcode_type, 16#0F#),
      1171 => to_slv(opcode_type, 16#0B#),
      1172 => to_slv(opcode_type, 16#09#),
      1173 => to_slv(opcode_type, 16#0B#),
      1174 => to_slv(opcode_type, 16#0C#),
      1175 => to_slv(opcode_type, 16#09#),
      1176 => to_slv(opcode_type, 16#09#),
      1177 => to_slv(opcode_type, 16#0D#),
      1178 => to_slv(opcode_type, 16#0F#),
      1179 => to_slv(opcode_type, 16#07#),
      1180 => to_slv(opcode_type, 16#0B#),
      1181 => to_slv(opcode_type, 16#0B#),
      1182 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#09#),
      1185 => to_slv(opcode_type, 16#09#),
      1186 => to_slv(opcode_type, 16#08#),
      1187 => to_slv(opcode_type, 16#04#),
      1188 => to_slv(opcode_type, 16#0F#),
      1189 => to_slv(opcode_type, 16#09#),
      1190 => to_slv(opcode_type, 16#0E#),
      1191 => to_slv(opcode_type, 16#0C#),
      1192 => to_slv(opcode_type, 16#06#),
      1193 => to_slv(opcode_type, 16#08#),
      1194 => to_slv(opcode_type, 16#10#),
      1195 => to_slv(opcode_type, 16#0B#),
      1196 => to_slv(opcode_type, 16#08#),
      1197 => to_slv(opcode_type, 16#0A#),
      1198 => to_slv(opcode_type, 16#0C#),
      1199 => to_slv(opcode_type, 16#09#),
      1200 => to_slv(opcode_type, 16#09#),
      1201 => to_slv(opcode_type, 16#08#),
      1202 => to_slv(opcode_type, 16#56#),
      1203 => to_slv(opcode_type, 16#10#),
      1204 => to_slv(opcode_type, 16#08#),
      1205 => to_slv(opcode_type, 16#0B#),
      1206 => to_slv(opcode_type, 16#11#),
      1207 => to_slv(opcode_type, 16#07#),
      1208 => to_slv(opcode_type, 16#09#),
      1209 => to_slv(opcode_type, 16#0C#),
      1210 => to_slv(opcode_type, 16#81#),
      1211 => to_slv(opcode_type, 16#07#),
      1212 => to_slv(opcode_type, 16#0E#),
      1213 => to_slv(opcode_type, 16#0C#),
      1214 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#07#),
      1217 => to_slv(opcode_type, 16#06#),
      1218 => to_slv(opcode_type, 16#06#),
      1219 => to_slv(opcode_type, 16#09#),
      1220 => to_slv(opcode_type, 16#0A#),
      1221 => to_slv(opcode_type, 16#DF#),
      1222 => to_slv(opcode_type, 16#06#),
      1223 => to_slv(opcode_type, 16#0A#),
      1224 => to_slv(opcode_type, 16#0B#),
      1225 => to_slv(opcode_type, 16#08#),
      1226 => to_slv(opcode_type, 16#08#),
      1227 => to_slv(opcode_type, 16#0A#),
      1228 => to_slv(opcode_type, 16#0A#),
      1229 => to_slv(opcode_type, 16#01#),
      1230 => to_slv(opcode_type, 16#0D#),
      1231 => to_slv(opcode_type, 16#08#),
      1232 => to_slv(opcode_type, 16#09#),
      1233 => to_slv(opcode_type, 16#08#),
      1234 => to_slv(opcode_type, 16#0E#),
      1235 => to_slv(opcode_type, 16#0E#),
      1236 => to_slv(opcode_type, 16#07#),
      1237 => to_slv(opcode_type, 16#0F#),
      1238 => to_slv(opcode_type, 16#0A#),
      1239 => to_slv(opcode_type, 16#06#),
      1240 => to_slv(opcode_type, 16#09#),
      1241 => to_slv(opcode_type, 16#0C#),
      1242 => to_slv(opcode_type, 16#0B#),
      1243 => to_slv(opcode_type, 16#08#),
      1244 => to_slv(opcode_type, 16#0B#),
      1245 => to_slv(opcode_type, 16#0C#),
      1246 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#06#),
      1249 => to_slv(opcode_type, 16#07#),
      1250 => to_slv(opcode_type, 16#07#),
      1251 => to_slv(opcode_type, 16#09#),
      1252 => to_slv(opcode_type, 16#0C#),
      1253 => to_slv(opcode_type, 16#0B#),
      1254 => to_slv(opcode_type, 16#07#),
      1255 => to_slv(opcode_type, 16#11#),
      1256 => to_slv(opcode_type, 16#11#),
      1257 => to_slv(opcode_type, 16#08#),
      1258 => to_slv(opcode_type, 16#01#),
      1259 => to_slv(opcode_type, 16#0A#),
      1260 => to_slv(opcode_type, 16#07#),
      1261 => to_slv(opcode_type, 16#10#),
      1262 => to_slv(opcode_type, 16#0C#),
      1263 => to_slv(opcode_type, 16#09#),
      1264 => to_slv(opcode_type, 16#08#),
      1265 => to_slv(opcode_type, 16#08#),
      1266 => to_slv(opcode_type, 16#0D#),
      1267 => to_slv(opcode_type, 16#10#),
      1268 => to_slv(opcode_type, 16#06#),
      1269 => to_slv(opcode_type, 16#10#),
      1270 => to_slv(opcode_type, 16#0F#),
      1271 => to_slv(opcode_type, 16#07#),
      1272 => to_slv(opcode_type, 16#08#),
      1273 => to_slv(opcode_type, 16#0D#),
      1274 => to_slv(opcode_type, 16#10#),
      1275 => to_slv(opcode_type, 16#09#),
      1276 => to_slv(opcode_type, 16#0D#),
      1277 => to_slv(opcode_type, 16#0C#),
      1278 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#06#),
      1281 => to_slv(opcode_type, 16#09#),
      1282 => to_slv(opcode_type, 16#09#),
      1283 => to_slv(opcode_type, 16#09#),
      1284 => to_slv(opcode_type, 16#0B#),
      1285 => to_slv(opcode_type, 16#10#),
      1286 => to_slv(opcode_type, 16#01#),
      1287 => to_slv(opcode_type, 16#0A#),
      1288 => to_slv(opcode_type, 16#06#),
      1289 => to_slv(opcode_type, 16#07#),
      1290 => to_slv(opcode_type, 16#0B#),
      1291 => to_slv(opcode_type, 16#0D#),
      1292 => to_slv(opcode_type, 16#09#),
      1293 => to_slv(opcode_type, 16#0B#),
      1294 => to_slv(opcode_type, 16#11#),
      1295 => to_slv(opcode_type, 16#08#),
      1296 => to_slv(opcode_type, 16#07#),
      1297 => to_slv(opcode_type, 16#07#),
      1298 => to_slv(opcode_type, 16#0B#),
      1299 => to_slv(opcode_type, 16#0E#),
      1300 => to_slv(opcode_type, 16#06#),
      1301 => to_slv(opcode_type, 16#52#),
      1302 => to_slv(opcode_type, 16#0E#),
      1303 => to_slv(opcode_type, 16#06#),
      1304 => to_slv(opcode_type, 16#07#),
      1305 => to_slv(opcode_type, 16#0F#),
      1306 => to_slv(opcode_type, 16#0C#),
      1307 => to_slv(opcode_type, 16#06#),
      1308 => to_slv(opcode_type, 16#0D#),
      1309 => to_slv(opcode_type, 16#11#),
      1310 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#07#),
      1313 => to_slv(opcode_type, 16#09#),
      1314 => to_slv(opcode_type, 16#07#),
      1315 => to_slv(opcode_type, 16#08#),
      1316 => to_slv(opcode_type, 16#0C#),
      1317 => to_slv(opcode_type, 16#AF#),
      1318 => to_slv(opcode_type, 16#07#),
      1319 => to_slv(opcode_type, 16#11#),
      1320 => to_slv(opcode_type, 16#0E#),
      1321 => to_slv(opcode_type, 16#08#),
      1322 => to_slv(opcode_type, 16#04#),
      1323 => to_slv(opcode_type, 16#0B#),
      1324 => to_slv(opcode_type, 16#07#),
      1325 => to_slv(opcode_type, 16#0F#),
      1326 => to_slv(opcode_type, 16#0F#),
      1327 => to_slv(opcode_type, 16#08#),
      1328 => to_slv(opcode_type, 16#08#),
      1329 => to_slv(opcode_type, 16#07#),
      1330 => to_slv(opcode_type, 16#0E#),
      1331 => to_slv(opcode_type, 16#0C#),
      1332 => to_slv(opcode_type, 16#09#),
      1333 => to_slv(opcode_type, 16#0A#),
      1334 => to_slv(opcode_type, 16#0C#),
      1335 => to_slv(opcode_type, 16#06#),
      1336 => to_slv(opcode_type, 16#09#),
      1337 => to_slv(opcode_type, 16#10#),
      1338 => to_slv(opcode_type, 16#0D#),
      1339 => to_slv(opcode_type, 16#09#),
      1340 => to_slv(opcode_type, 16#0E#),
      1341 => to_slv(opcode_type, 16#0A#),
      1342 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#09#),
      1345 => to_slv(opcode_type, 16#09#),
      1346 => to_slv(opcode_type, 16#08#),
      1347 => to_slv(opcode_type, 16#06#),
      1348 => to_slv(opcode_type, 16#0D#),
      1349 => to_slv(opcode_type, 16#10#),
      1350 => to_slv(opcode_type, 16#05#),
      1351 => to_slv(opcode_type, 16#5C#),
      1352 => to_slv(opcode_type, 16#09#),
      1353 => to_slv(opcode_type, 16#08#),
      1354 => to_slv(opcode_type, 16#0B#),
      1355 => to_slv(opcode_type, 16#0F#),
      1356 => to_slv(opcode_type, 16#09#),
      1357 => to_slv(opcode_type, 16#0C#),
      1358 => to_slv(opcode_type, 16#8A#),
      1359 => to_slv(opcode_type, 16#09#),
      1360 => to_slv(opcode_type, 16#09#),
      1361 => to_slv(opcode_type, 16#09#),
      1362 => to_slv(opcode_type, 16#0F#),
      1363 => to_slv(opcode_type, 16#11#),
      1364 => to_slv(opcode_type, 16#09#),
      1365 => to_slv(opcode_type, 16#0B#),
      1366 => to_slv(opcode_type, 16#0C#),
      1367 => to_slv(opcode_type, 16#09#),
      1368 => to_slv(opcode_type, 16#09#),
      1369 => to_slv(opcode_type, 16#10#),
      1370 => to_slv(opcode_type, 16#0A#),
      1371 => to_slv(opcode_type, 16#06#),
      1372 => to_slv(opcode_type, 16#0A#),
      1373 => to_slv(opcode_type, 16#0B#),
      1374 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#06#),
      1377 => to_slv(opcode_type, 16#06#),
      1378 => to_slv(opcode_type, 16#06#),
      1379 => to_slv(opcode_type, 16#09#),
      1380 => to_slv(opcode_type, 16#0D#),
      1381 => to_slv(opcode_type, 16#B8#),
      1382 => to_slv(opcode_type, 16#04#),
      1383 => to_slv(opcode_type, 16#0D#),
      1384 => to_slv(opcode_type, 16#08#),
      1385 => to_slv(opcode_type, 16#09#),
      1386 => to_slv(opcode_type, 16#0B#),
      1387 => to_slv(opcode_type, 16#3D#),
      1388 => to_slv(opcode_type, 16#09#),
      1389 => to_slv(opcode_type, 16#10#),
      1390 => to_slv(opcode_type, 16#0B#),
      1391 => to_slv(opcode_type, 16#07#),
      1392 => to_slv(opcode_type, 16#09#),
      1393 => to_slv(opcode_type, 16#07#),
      1394 => to_slv(opcode_type, 16#0A#),
      1395 => to_slv(opcode_type, 16#34#),
      1396 => to_slv(opcode_type, 16#06#),
      1397 => to_slv(opcode_type, 16#0F#),
      1398 => to_slv(opcode_type, 16#0D#),
      1399 => to_slv(opcode_type, 16#07#),
      1400 => to_slv(opcode_type, 16#08#),
      1401 => to_slv(opcode_type, 16#0B#),
      1402 => to_slv(opcode_type, 16#0B#),
      1403 => to_slv(opcode_type, 16#09#),
      1404 => to_slv(opcode_type, 16#10#),
      1405 => to_slv(opcode_type, 16#11#),
      1406 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#06#),
      1409 => to_slv(opcode_type, 16#07#),
      1410 => to_slv(opcode_type, 16#06#),
      1411 => to_slv(opcode_type, 16#07#),
      1412 => to_slv(opcode_type, 16#0A#),
      1413 => to_slv(opcode_type, 16#0D#),
      1414 => to_slv(opcode_type, 16#02#),
      1415 => to_slv(opcode_type, 16#11#),
      1416 => to_slv(opcode_type, 16#09#),
      1417 => to_slv(opcode_type, 16#08#),
      1418 => to_slv(opcode_type, 16#0A#),
      1419 => to_slv(opcode_type, 16#6A#),
      1420 => to_slv(opcode_type, 16#08#),
      1421 => to_slv(opcode_type, 16#0A#),
      1422 => to_slv(opcode_type, 16#0D#),
      1423 => to_slv(opcode_type, 16#06#),
      1424 => to_slv(opcode_type, 16#07#),
      1425 => to_slv(opcode_type, 16#09#),
      1426 => to_slv(opcode_type, 16#0C#),
      1427 => to_slv(opcode_type, 16#11#),
      1428 => to_slv(opcode_type, 16#08#),
      1429 => to_slv(opcode_type, 16#0C#),
      1430 => to_slv(opcode_type, 16#7A#),
      1431 => to_slv(opcode_type, 16#08#),
      1432 => to_slv(opcode_type, 16#09#),
      1433 => to_slv(opcode_type, 16#10#),
      1434 => to_slv(opcode_type, 16#0A#),
      1435 => to_slv(opcode_type, 16#09#),
      1436 => to_slv(opcode_type, 16#0F#),
      1437 => to_slv(opcode_type, 16#0C#),
      1438 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#08#),
      1441 => to_slv(opcode_type, 16#08#),
      1442 => to_slv(opcode_type, 16#08#),
      1443 => to_slv(opcode_type, 16#05#),
      1444 => to_slv(opcode_type, 16#0E#),
      1445 => to_slv(opcode_type, 16#06#),
      1446 => to_slv(opcode_type, 16#0A#),
      1447 => to_slv(opcode_type, 16#EC#),
      1448 => to_slv(opcode_type, 16#06#),
      1449 => to_slv(opcode_type, 16#08#),
      1450 => to_slv(opcode_type, 16#0A#),
      1451 => to_slv(opcode_type, 16#0F#),
      1452 => to_slv(opcode_type, 16#06#),
      1453 => to_slv(opcode_type, 16#0F#),
      1454 => to_slv(opcode_type, 16#0A#),
      1455 => to_slv(opcode_type, 16#08#),
      1456 => to_slv(opcode_type, 16#06#),
      1457 => to_slv(opcode_type, 16#09#),
      1458 => to_slv(opcode_type, 16#0C#),
      1459 => to_slv(opcode_type, 16#D8#),
      1460 => to_slv(opcode_type, 16#07#),
      1461 => to_slv(opcode_type, 16#0F#),
      1462 => to_slv(opcode_type, 16#0A#),
      1463 => to_slv(opcode_type, 16#06#),
      1464 => to_slv(opcode_type, 16#09#),
      1465 => to_slv(opcode_type, 16#10#),
      1466 => to_slv(opcode_type, 16#11#),
      1467 => to_slv(opcode_type, 16#07#),
      1468 => to_slv(opcode_type, 16#0F#),
      1469 => to_slv(opcode_type, 16#0A#),
      1470 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#07#),
      1473 => to_slv(opcode_type, 16#09#),
      1474 => to_slv(opcode_type, 16#07#),
      1475 => to_slv(opcode_type, 16#06#),
      1476 => to_slv(opcode_type, 16#0F#),
      1477 => to_slv(opcode_type, 16#0A#),
      1478 => to_slv(opcode_type, 16#02#),
      1479 => to_slv(opcode_type, 16#8E#),
      1480 => to_slv(opcode_type, 16#07#),
      1481 => to_slv(opcode_type, 16#08#),
      1482 => to_slv(opcode_type, 16#0C#),
      1483 => to_slv(opcode_type, 16#10#),
      1484 => to_slv(opcode_type, 16#06#),
      1485 => to_slv(opcode_type, 16#10#),
      1486 => to_slv(opcode_type, 16#FC#),
      1487 => to_slv(opcode_type, 16#07#),
      1488 => to_slv(opcode_type, 16#06#),
      1489 => to_slv(opcode_type, 16#08#),
      1490 => to_slv(opcode_type, 16#11#),
      1491 => to_slv(opcode_type, 16#10#),
      1492 => to_slv(opcode_type, 16#06#),
      1493 => to_slv(opcode_type, 16#0E#),
      1494 => to_slv(opcode_type, 16#AA#),
      1495 => to_slv(opcode_type, 16#07#),
      1496 => to_slv(opcode_type, 16#06#),
      1497 => to_slv(opcode_type, 16#0C#),
      1498 => to_slv(opcode_type, 16#0B#),
      1499 => to_slv(opcode_type, 16#08#),
      1500 => to_slv(opcode_type, 16#0B#),
      1501 => to_slv(opcode_type, 16#12#),
      1502 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#06#),
      1505 => to_slv(opcode_type, 16#06#),
      1506 => to_slv(opcode_type, 16#07#),
      1507 => to_slv(opcode_type, 16#06#),
      1508 => to_slv(opcode_type, 16#11#),
      1509 => to_slv(opcode_type, 16#10#),
      1510 => to_slv(opcode_type, 16#04#),
      1511 => to_slv(opcode_type, 16#0F#),
      1512 => to_slv(opcode_type, 16#09#),
      1513 => to_slv(opcode_type, 16#08#),
      1514 => to_slv(opcode_type, 16#D1#),
      1515 => to_slv(opcode_type, 16#11#),
      1516 => to_slv(opcode_type, 16#07#),
      1517 => to_slv(opcode_type, 16#0A#),
      1518 => to_slv(opcode_type, 16#11#),
      1519 => to_slv(opcode_type, 16#06#),
      1520 => to_slv(opcode_type, 16#07#),
      1521 => to_slv(opcode_type, 16#06#),
      1522 => to_slv(opcode_type, 16#11#),
      1523 => to_slv(opcode_type, 16#0A#),
      1524 => to_slv(opcode_type, 16#06#),
      1525 => to_slv(opcode_type, 16#0B#),
      1526 => to_slv(opcode_type, 16#0D#),
      1527 => to_slv(opcode_type, 16#07#),
      1528 => to_slv(opcode_type, 16#08#),
      1529 => to_slv(opcode_type, 16#D9#),
      1530 => to_slv(opcode_type, 16#0E#),
      1531 => to_slv(opcode_type, 16#08#),
      1532 => to_slv(opcode_type, 16#0A#),
      1533 => to_slv(opcode_type, 16#10#),
      1534 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#07#),
      1537 => to_slv(opcode_type, 16#08#),
      1538 => to_slv(opcode_type, 16#08#),
      1539 => to_slv(opcode_type, 16#05#),
      1540 => to_slv(opcode_type, 16#0D#),
      1541 => to_slv(opcode_type, 16#09#),
      1542 => to_slv(opcode_type, 16#0A#),
      1543 => to_slv(opcode_type, 16#0A#),
      1544 => to_slv(opcode_type, 16#09#),
      1545 => to_slv(opcode_type, 16#07#),
      1546 => to_slv(opcode_type, 16#10#),
      1547 => to_slv(opcode_type, 16#11#),
      1548 => to_slv(opcode_type, 16#09#),
      1549 => to_slv(opcode_type, 16#0C#),
      1550 => to_slv(opcode_type, 16#0E#),
      1551 => to_slv(opcode_type, 16#06#),
      1552 => to_slv(opcode_type, 16#09#),
      1553 => to_slv(opcode_type, 16#07#),
      1554 => to_slv(opcode_type, 16#0F#),
      1555 => to_slv(opcode_type, 16#0E#),
      1556 => to_slv(opcode_type, 16#09#),
      1557 => to_slv(opcode_type, 16#0F#),
      1558 => to_slv(opcode_type, 16#0E#),
      1559 => to_slv(opcode_type, 16#07#),
      1560 => to_slv(opcode_type, 16#07#),
      1561 => to_slv(opcode_type, 16#0A#),
      1562 => to_slv(opcode_type, 16#0A#),
      1563 => to_slv(opcode_type, 16#09#),
      1564 => to_slv(opcode_type, 16#11#),
      1565 => to_slv(opcode_type, 16#0A#),
      1566 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#07#),
      1569 => to_slv(opcode_type, 16#06#),
      1570 => to_slv(opcode_type, 16#07#),
      1571 => to_slv(opcode_type, 16#09#),
      1572 => to_slv(opcode_type, 16#0F#),
      1573 => to_slv(opcode_type, 16#0C#),
      1574 => to_slv(opcode_type, 16#06#),
      1575 => to_slv(opcode_type, 16#0E#),
      1576 => to_slv(opcode_type, 16#10#),
      1577 => to_slv(opcode_type, 16#07#),
      1578 => to_slv(opcode_type, 16#01#),
      1579 => to_slv(opcode_type, 16#0F#),
      1580 => to_slv(opcode_type, 16#09#),
      1581 => to_slv(opcode_type, 16#0C#),
      1582 => to_slv(opcode_type, 16#0B#),
      1583 => to_slv(opcode_type, 16#08#),
      1584 => to_slv(opcode_type, 16#09#),
      1585 => to_slv(opcode_type, 16#06#),
      1586 => to_slv(opcode_type, 16#DD#),
      1587 => to_slv(opcode_type, 16#0F#),
      1588 => to_slv(opcode_type, 16#08#),
      1589 => to_slv(opcode_type, 16#96#),
      1590 => to_slv(opcode_type, 16#0B#),
      1591 => to_slv(opcode_type, 16#09#),
      1592 => to_slv(opcode_type, 16#06#),
      1593 => to_slv(opcode_type, 16#0F#),
      1594 => to_slv(opcode_type, 16#0C#),
      1595 => to_slv(opcode_type, 16#08#),
      1596 => to_slv(opcode_type, 16#0C#),
      1597 => to_slv(opcode_type, 16#0A#),
      1598 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#07#),
      1602 => to_slv(opcode_type, 16#07#),
      1603 => to_slv(opcode_type, 16#05#),
      1604 => to_slv(opcode_type, 16#0E#),
      1605 => to_slv(opcode_type, 16#09#),
      1606 => to_slv(opcode_type, 16#0F#),
      1607 => to_slv(opcode_type, 16#EA#),
      1608 => to_slv(opcode_type, 16#06#),
      1609 => to_slv(opcode_type, 16#06#),
      1610 => to_slv(opcode_type, 16#10#),
      1611 => to_slv(opcode_type, 16#0F#),
      1612 => to_slv(opcode_type, 16#07#),
      1613 => to_slv(opcode_type, 16#0E#),
      1614 => to_slv(opcode_type, 16#0D#),
      1615 => to_slv(opcode_type, 16#06#),
      1616 => to_slv(opcode_type, 16#08#),
      1617 => to_slv(opcode_type, 16#09#),
      1618 => to_slv(opcode_type, 16#0F#),
      1619 => to_slv(opcode_type, 16#0B#),
      1620 => to_slv(opcode_type, 16#09#),
      1621 => to_slv(opcode_type, 16#10#),
      1622 => to_slv(opcode_type, 16#10#),
      1623 => to_slv(opcode_type, 16#07#),
      1624 => to_slv(opcode_type, 16#07#),
      1625 => to_slv(opcode_type, 16#10#),
      1626 => to_slv(opcode_type, 16#11#),
      1627 => to_slv(opcode_type, 16#07#),
      1628 => to_slv(opcode_type, 16#0B#),
      1629 => to_slv(opcode_type, 16#0A#),
      1630 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#09#),
      1633 => to_slv(opcode_type, 16#08#),
      1634 => to_slv(opcode_type, 16#08#),
      1635 => to_slv(opcode_type, 16#07#),
      1636 => to_slv(opcode_type, 16#0F#),
      1637 => to_slv(opcode_type, 16#F5#),
      1638 => to_slv(opcode_type, 16#08#),
      1639 => to_slv(opcode_type, 16#10#),
      1640 => to_slv(opcode_type, 16#0B#),
      1641 => to_slv(opcode_type, 16#08#),
      1642 => to_slv(opcode_type, 16#03#),
      1643 => to_slv(opcode_type, 16#0C#),
      1644 => to_slv(opcode_type, 16#06#),
      1645 => to_slv(opcode_type, 16#0D#),
      1646 => to_slv(opcode_type, 16#0B#),
      1647 => to_slv(opcode_type, 16#08#),
      1648 => to_slv(opcode_type, 16#08#),
      1649 => to_slv(opcode_type, 16#09#),
      1650 => to_slv(opcode_type, 16#0E#),
      1651 => to_slv(opcode_type, 16#0E#),
      1652 => to_slv(opcode_type, 16#09#),
      1653 => to_slv(opcode_type, 16#7E#),
      1654 => to_slv(opcode_type, 16#0D#),
      1655 => to_slv(opcode_type, 16#09#),
      1656 => to_slv(opcode_type, 16#07#),
      1657 => to_slv(opcode_type, 16#0A#),
      1658 => to_slv(opcode_type, 16#0A#),
      1659 => to_slv(opcode_type, 16#06#),
      1660 => to_slv(opcode_type, 16#0E#),
      1661 => to_slv(opcode_type, 16#0D#),
      1662 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#09#),
      1665 => to_slv(opcode_type, 16#08#),
      1666 => to_slv(opcode_type, 16#07#),
      1667 => to_slv(opcode_type, 16#04#),
      1668 => to_slv(opcode_type, 16#0E#),
      1669 => to_slv(opcode_type, 16#09#),
      1670 => to_slv(opcode_type, 16#0B#),
      1671 => to_slv(opcode_type, 16#0D#),
      1672 => to_slv(opcode_type, 16#07#),
      1673 => to_slv(opcode_type, 16#09#),
      1674 => to_slv(opcode_type, 16#0F#),
      1675 => to_slv(opcode_type, 16#0C#),
      1676 => to_slv(opcode_type, 16#09#),
      1677 => to_slv(opcode_type, 16#0D#),
      1678 => to_slv(opcode_type, 16#10#),
      1679 => to_slv(opcode_type, 16#07#),
      1680 => to_slv(opcode_type, 16#08#),
      1681 => to_slv(opcode_type, 16#06#),
      1682 => to_slv(opcode_type, 16#0E#),
      1683 => to_slv(opcode_type, 16#10#),
      1684 => to_slv(opcode_type, 16#08#),
      1685 => to_slv(opcode_type, 16#0D#),
      1686 => to_slv(opcode_type, 16#0C#),
      1687 => to_slv(opcode_type, 16#09#),
      1688 => to_slv(opcode_type, 16#06#),
      1689 => to_slv(opcode_type, 16#DC#),
      1690 => to_slv(opcode_type, 16#6A#),
      1691 => to_slv(opcode_type, 16#08#),
      1692 => to_slv(opcode_type, 16#0F#),
      1693 => to_slv(opcode_type, 16#11#),
      1694 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#09#),
      1697 => to_slv(opcode_type, 16#09#),
      1698 => to_slv(opcode_type, 16#06#),
      1699 => to_slv(opcode_type, 16#01#),
      1700 => to_slv(opcode_type, 16#0A#),
      1701 => to_slv(opcode_type, 16#08#),
      1702 => to_slv(opcode_type, 16#0C#),
      1703 => to_slv(opcode_type, 16#11#),
      1704 => to_slv(opcode_type, 16#08#),
      1705 => to_slv(opcode_type, 16#09#),
      1706 => to_slv(opcode_type, 16#F6#),
      1707 => to_slv(opcode_type, 16#0B#),
      1708 => to_slv(opcode_type, 16#07#),
      1709 => to_slv(opcode_type, 16#11#),
      1710 => to_slv(opcode_type, 16#10#),
      1711 => to_slv(opcode_type, 16#07#),
      1712 => to_slv(opcode_type, 16#08#),
      1713 => to_slv(opcode_type, 16#09#),
      1714 => to_slv(opcode_type, 16#0D#),
      1715 => to_slv(opcode_type, 16#0D#),
      1716 => to_slv(opcode_type, 16#06#),
      1717 => to_slv(opcode_type, 16#0C#),
      1718 => to_slv(opcode_type, 16#10#),
      1719 => to_slv(opcode_type, 16#08#),
      1720 => to_slv(opcode_type, 16#06#),
      1721 => to_slv(opcode_type, 16#0D#),
      1722 => to_slv(opcode_type, 16#0D#),
      1723 => to_slv(opcode_type, 16#09#),
      1724 => to_slv(opcode_type, 16#10#),
      1725 => to_slv(opcode_type, 16#0A#),
      1726 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#07#),
      1729 => to_slv(opcode_type, 16#09#),
      1730 => to_slv(opcode_type, 16#08#),
      1731 => to_slv(opcode_type, 16#05#),
      1732 => to_slv(opcode_type, 16#0C#),
      1733 => to_slv(opcode_type, 16#06#),
      1734 => to_slv(opcode_type, 16#0C#),
      1735 => to_slv(opcode_type, 16#11#),
      1736 => to_slv(opcode_type, 16#07#),
      1737 => to_slv(opcode_type, 16#07#),
      1738 => to_slv(opcode_type, 16#10#),
      1739 => to_slv(opcode_type, 16#11#),
      1740 => to_slv(opcode_type, 16#09#),
      1741 => to_slv(opcode_type, 16#10#),
      1742 => to_slv(opcode_type, 16#0B#),
      1743 => to_slv(opcode_type, 16#08#),
      1744 => to_slv(opcode_type, 16#07#),
      1745 => to_slv(opcode_type, 16#08#),
      1746 => to_slv(opcode_type, 16#0B#),
      1747 => to_slv(opcode_type, 16#C7#),
      1748 => to_slv(opcode_type, 16#06#),
      1749 => to_slv(opcode_type, 16#0A#),
      1750 => to_slv(opcode_type, 16#0A#),
      1751 => to_slv(opcode_type, 16#09#),
      1752 => to_slv(opcode_type, 16#09#),
      1753 => to_slv(opcode_type, 16#0A#),
      1754 => to_slv(opcode_type, 16#0A#),
      1755 => to_slv(opcode_type, 16#06#),
      1756 => to_slv(opcode_type, 16#89#),
      1757 => to_slv(opcode_type, 16#0E#),
      1758 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#06#),
      1761 => to_slv(opcode_type, 16#08#),
      1762 => to_slv(opcode_type, 16#06#),
      1763 => to_slv(opcode_type, 16#02#),
      1764 => to_slv(opcode_type, 16#0D#),
      1765 => to_slv(opcode_type, 16#09#),
      1766 => to_slv(opcode_type, 16#10#),
      1767 => to_slv(opcode_type, 16#0A#),
      1768 => to_slv(opcode_type, 16#06#),
      1769 => to_slv(opcode_type, 16#08#),
      1770 => to_slv(opcode_type, 16#D0#),
      1771 => to_slv(opcode_type, 16#0C#),
      1772 => to_slv(opcode_type, 16#08#),
      1773 => to_slv(opcode_type, 16#0A#),
      1774 => to_slv(opcode_type, 16#0F#),
      1775 => to_slv(opcode_type, 16#09#),
      1776 => to_slv(opcode_type, 16#09#),
      1777 => to_slv(opcode_type, 16#08#),
      1778 => to_slv(opcode_type, 16#11#),
      1779 => to_slv(opcode_type, 16#0B#),
      1780 => to_slv(opcode_type, 16#09#),
      1781 => to_slv(opcode_type, 16#11#),
      1782 => to_slv(opcode_type, 16#0C#),
      1783 => to_slv(opcode_type, 16#07#),
      1784 => to_slv(opcode_type, 16#09#),
      1785 => to_slv(opcode_type, 16#0C#),
      1786 => to_slv(opcode_type, 16#0A#),
      1787 => to_slv(opcode_type, 16#09#),
      1788 => to_slv(opcode_type, 16#6A#),
      1789 => to_slv(opcode_type, 16#0C#),
      1790 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#08#),
      1793 => to_slv(opcode_type, 16#09#),
      1794 => to_slv(opcode_type, 16#09#),
      1795 => to_slv(opcode_type, 16#07#),
      1796 => to_slv(opcode_type, 16#0E#),
      1797 => to_slv(opcode_type, 16#11#),
      1798 => to_slv(opcode_type, 16#06#),
      1799 => to_slv(opcode_type, 16#0F#),
      1800 => to_slv(opcode_type, 16#0D#),
      1801 => to_slv(opcode_type, 16#08#),
      1802 => to_slv(opcode_type, 16#05#),
      1803 => to_slv(opcode_type, 16#10#),
      1804 => to_slv(opcode_type, 16#08#),
      1805 => to_slv(opcode_type, 16#0D#),
      1806 => to_slv(opcode_type, 16#11#),
      1807 => to_slv(opcode_type, 16#08#),
      1808 => to_slv(opcode_type, 16#09#),
      1809 => to_slv(opcode_type, 16#06#),
      1810 => to_slv(opcode_type, 16#0C#),
      1811 => to_slv(opcode_type, 16#0D#),
      1812 => to_slv(opcode_type, 16#09#),
      1813 => to_slv(opcode_type, 16#0A#),
      1814 => to_slv(opcode_type, 16#0D#),
      1815 => to_slv(opcode_type, 16#07#),
      1816 => to_slv(opcode_type, 16#08#),
      1817 => to_slv(opcode_type, 16#10#),
      1818 => to_slv(opcode_type, 16#10#),
      1819 => to_slv(opcode_type, 16#06#),
      1820 => to_slv(opcode_type, 16#0F#),
      1821 => to_slv(opcode_type, 16#0E#),
      1822 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#06#),
      1825 => to_slv(opcode_type, 16#08#),
      1826 => to_slv(opcode_type, 16#06#),
      1827 => to_slv(opcode_type, 16#07#),
      1828 => to_slv(opcode_type, 16#0D#),
      1829 => to_slv(opcode_type, 16#11#),
      1830 => to_slv(opcode_type, 16#08#),
      1831 => to_slv(opcode_type, 16#0F#),
      1832 => to_slv(opcode_type, 16#0E#),
      1833 => to_slv(opcode_type, 16#08#),
      1834 => to_slv(opcode_type, 16#01#),
      1835 => to_slv(opcode_type, 16#0E#),
      1836 => to_slv(opcode_type, 16#06#),
      1837 => to_slv(opcode_type, 16#0D#),
      1838 => to_slv(opcode_type, 16#0A#),
      1839 => to_slv(opcode_type, 16#06#),
      1840 => to_slv(opcode_type, 16#06#),
      1841 => to_slv(opcode_type, 16#06#),
      1842 => to_slv(opcode_type, 16#DF#),
      1843 => to_slv(opcode_type, 16#0D#),
      1844 => to_slv(opcode_type, 16#08#),
      1845 => to_slv(opcode_type, 16#11#),
      1846 => to_slv(opcode_type, 16#0D#),
      1847 => to_slv(opcode_type, 16#08#),
      1848 => to_slv(opcode_type, 16#09#),
      1849 => to_slv(opcode_type, 16#0F#),
      1850 => to_slv(opcode_type, 16#0B#),
      1851 => to_slv(opcode_type, 16#08#),
      1852 => to_slv(opcode_type, 16#0D#),
      1853 => to_slv(opcode_type, 16#C1#),
      1854 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#09#),
      1857 => to_slv(opcode_type, 16#07#),
      1858 => to_slv(opcode_type, 16#09#),
      1859 => to_slv(opcode_type, 16#07#),
      1860 => to_slv(opcode_type, 16#0C#),
      1861 => to_slv(opcode_type, 16#0A#),
      1862 => to_slv(opcode_type, 16#04#),
      1863 => to_slv(opcode_type, 16#4A#),
      1864 => to_slv(opcode_type, 16#06#),
      1865 => to_slv(opcode_type, 16#09#),
      1866 => to_slv(opcode_type, 16#0A#),
      1867 => to_slv(opcode_type, 16#0F#),
      1868 => to_slv(opcode_type, 16#09#),
      1869 => to_slv(opcode_type, 16#0C#),
      1870 => to_slv(opcode_type, 16#0C#),
      1871 => to_slv(opcode_type, 16#08#),
      1872 => to_slv(opcode_type, 16#07#),
      1873 => to_slv(opcode_type, 16#09#),
      1874 => to_slv(opcode_type, 16#0C#),
      1875 => to_slv(opcode_type, 16#10#),
      1876 => to_slv(opcode_type, 16#06#),
      1877 => to_slv(opcode_type, 16#0E#),
      1878 => to_slv(opcode_type, 16#10#),
      1879 => to_slv(opcode_type, 16#08#),
      1880 => to_slv(opcode_type, 16#08#),
      1881 => to_slv(opcode_type, 16#0E#),
      1882 => to_slv(opcode_type, 16#0D#),
      1883 => to_slv(opcode_type, 16#07#),
      1884 => to_slv(opcode_type, 16#10#),
      1885 => to_slv(opcode_type, 16#0A#),
      1886 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#08#),
      1890 => to_slv(opcode_type, 16#06#),
      1891 => to_slv(opcode_type, 16#01#),
      1892 => to_slv(opcode_type, 16#0E#),
      1893 => to_slv(opcode_type, 16#06#),
      1894 => to_slv(opcode_type, 16#0A#),
      1895 => to_slv(opcode_type, 16#0D#),
      1896 => to_slv(opcode_type, 16#07#),
      1897 => to_slv(opcode_type, 16#06#),
      1898 => to_slv(opcode_type, 16#0C#),
      1899 => to_slv(opcode_type, 16#0F#),
      1900 => to_slv(opcode_type, 16#08#),
      1901 => to_slv(opcode_type, 16#0C#),
      1902 => to_slv(opcode_type, 16#0B#),
      1903 => to_slv(opcode_type, 16#08#),
      1904 => to_slv(opcode_type, 16#08#),
      1905 => to_slv(opcode_type, 16#06#),
      1906 => to_slv(opcode_type, 16#0F#),
      1907 => to_slv(opcode_type, 16#0E#),
      1908 => to_slv(opcode_type, 16#08#),
      1909 => to_slv(opcode_type, 16#10#),
      1910 => to_slv(opcode_type, 16#11#),
      1911 => to_slv(opcode_type, 16#06#),
      1912 => to_slv(opcode_type, 16#06#),
      1913 => to_slv(opcode_type, 16#E4#),
      1914 => to_slv(opcode_type, 16#0C#),
      1915 => to_slv(opcode_type, 16#06#),
      1916 => to_slv(opcode_type, 16#0B#),
      1917 => to_slv(opcode_type, 16#10#),
      1918 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#06#),
      1921 => to_slv(opcode_type, 16#09#),
      1922 => to_slv(opcode_type, 16#09#),
      1923 => to_slv(opcode_type, 16#02#),
      1924 => to_slv(opcode_type, 16#0A#),
      1925 => to_slv(opcode_type, 16#07#),
      1926 => to_slv(opcode_type, 16#10#),
      1927 => to_slv(opcode_type, 16#0A#),
      1928 => to_slv(opcode_type, 16#06#),
      1929 => to_slv(opcode_type, 16#06#),
      1930 => to_slv(opcode_type, 16#1D#),
      1931 => to_slv(opcode_type, 16#0C#),
      1932 => to_slv(opcode_type, 16#08#),
      1933 => to_slv(opcode_type, 16#4B#),
      1934 => to_slv(opcode_type, 16#0C#),
      1935 => to_slv(opcode_type, 16#09#),
      1936 => to_slv(opcode_type, 16#09#),
      1937 => to_slv(opcode_type, 16#07#),
      1938 => to_slv(opcode_type, 16#0B#),
      1939 => to_slv(opcode_type, 16#0A#),
      1940 => to_slv(opcode_type, 16#09#),
      1941 => to_slv(opcode_type, 16#0E#),
      1942 => to_slv(opcode_type, 16#0E#),
      1943 => to_slv(opcode_type, 16#06#),
      1944 => to_slv(opcode_type, 16#09#),
      1945 => to_slv(opcode_type, 16#0B#),
      1946 => to_slv(opcode_type, 16#0A#),
      1947 => to_slv(opcode_type, 16#06#),
      1948 => to_slv(opcode_type, 16#0B#),
      1949 => to_slv(opcode_type, 16#0E#),
      1950 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#09#),
      1953 => to_slv(opcode_type, 16#06#),
      1954 => to_slv(opcode_type, 16#09#),
      1955 => to_slv(opcode_type, 16#05#),
      1956 => to_slv(opcode_type, 16#0A#),
      1957 => to_slv(opcode_type, 16#09#),
      1958 => to_slv(opcode_type, 16#11#),
      1959 => to_slv(opcode_type, 16#0D#),
      1960 => to_slv(opcode_type, 16#06#),
      1961 => to_slv(opcode_type, 16#08#),
      1962 => to_slv(opcode_type, 16#0D#),
      1963 => to_slv(opcode_type, 16#0C#),
      1964 => to_slv(opcode_type, 16#06#),
      1965 => to_slv(opcode_type, 16#11#),
      1966 => to_slv(opcode_type, 16#0A#),
      1967 => to_slv(opcode_type, 16#06#),
      1968 => to_slv(opcode_type, 16#06#),
      1969 => to_slv(opcode_type, 16#07#),
      1970 => to_slv(opcode_type, 16#11#),
      1971 => to_slv(opcode_type, 16#11#),
      1972 => to_slv(opcode_type, 16#06#),
      1973 => to_slv(opcode_type, 16#0E#),
      1974 => to_slv(opcode_type, 16#0E#),
      1975 => to_slv(opcode_type, 16#06#),
      1976 => to_slv(opcode_type, 16#08#),
      1977 => to_slv(opcode_type, 16#0F#),
      1978 => to_slv(opcode_type, 16#3E#),
      1979 => to_slv(opcode_type, 16#08#),
      1980 => to_slv(opcode_type, 16#35#),
      1981 => to_slv(opcode_type, 16#0D#),
      1982 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#07#),
      1985 => to_slv(opcode_type, 16#09#),
      1986 => to_slv(opcode_type, 16#07#),
      1987 => to_slv(opcode_type, 16#01#),
      1988 => to_slv(opcode_type, 16#10#),
      1989 => to_slv(opcode_type, 16#09#),
      1990 => to_slv(opcode_type, 16#0C#),
      1991 => to_slv(opcode_type, 16#0A#),
      1992 => to_slv(opcode_type, 16#06#),
      1993 => to_slv(opcode_type, 16#08#),
      1994 => to_slv(opcode_type, 16#AE#),
      1995 => to_slv(opcode_type, 16#11#),
      1996 => to_slv(opcode_type, 16#09#),
      1997 => to_slv(opcode_type, 16#0D#),
      1998 => to_slv(opcode_type, 16#0C#),
      1999 => to_slv(opcode_type, 16#08#),
      2000 => to_slv(opcode_type, 16#08#),
      2001 => to_slv(opcode_type, 16#08#),
      2002 => to_slv(opcode_type, 16#0D#),
      2003 => to_slv(opcode_type, 16#0D#),
      2004 => to_slv(opcode_type, 16#06#),
      2005 => to_slv(opcode_type, 16#0D#),
      2006 => to_slv(opcode_type, 16#0A#),
      2007 => to_slv(opcode_type, 16#06#),
      2008 => to_slv(opcode_type, 16#06#),
      2009 => to_slv(opcode_type, 16#F4#),
      2010 => to_slv(opcode_type, 16#0A#),
      2011 => to_slv(opcode_type, 16#06#),
      2012 => to_slv(opcode_type, 16#0E#),
      2013 => to_slv(opcode_type, 16#0B#),
      2014 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#07#),
      2017 => to_slv(opcode_type, 16#09#),
      2018 => to_slv(opcode_type, 16#07#),
      2019 => to_slv(opcode_type, 16#07#),
      2020 => to_slv(opcode_type, 16#0E#),
      2021 => to_slv(opcode_type, 16#10#),
      2022 => to_slv(opcode_type, 16#06#),
      2023 => to_slv(opcode_type, 16#0E#),
      2024 => to_slv(opcode_type, 16#0C#),
      2025 => to_slv(opcode_type, 16#09#),
      2026 => to_slv(opcode_type, 16#07#),
      2027 => to_slv(opcode_type, 16#0B#),
      2028 => to_slv(opcode_type, 16#10#),
      2029 => to_slv(opcode_type, 16#06#),
      2030 => to_slv(opcode_type, 16#0A#),
      2031 => to_slv(opcode_type, 16#10#),
      2032 => to_slv(opcode_type, 16#08#),
      2033 => to_slv(opcode_type, 16#08#),
      2034 => to_slv(opcode_type, 16#03#),
      2035 => to_slv(opcode_type, 16#11#),
      2036 => to_slv(opcode_type, 16#06#),
      2037 => to_slv(opcode_type, 16#11#),
      2038 => to_slv(opcode_type, 16#11#),
      2039 => to_slv(opcode_type, 16#09#),
      2040 => to_slv(opcode_type, 16#08#),
      2041 => to_slv(opcode_type, 16#0E#),
      2042 => to_slv(opcode_type, 16#11#),
      2043 => to_slv(opcode_type, 16#08#),
      2044 => to_slv(opcode_type, 16#0E#),
      2045 => to_slv(opcode_type, 16#0C#),
      2046 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#06#),
      2049 => to_slv(opcode_type, 16#07#),
      2050 => to_slv(opcode_type, 16#08#),
      2051 => to_slv(opcode_type, 16#01#),
      2052 => to_slv(opcode_type, 16#0C#),
      2053 => to_slv(opcode_type, 16#06#),
      2054 => to_slv(opcode_type, 16#0E#),
      2055 => to_slv(opcode_type, 16#10#),
      2056 => to_slv(opcode_type, 16#06#),
      2057 => to_slv(opcode_type, 16#07#),
      2058 => to_slv(opcode_type, 16#0A#),
      2059 => to_slv(opcode_type, 16#0A#),
      2060 => to_slv(opcode_type, 16#06#),
      2061 => to_slv(opcode_type, 16#10#),
      2062 => to_slv(opcode_type, 16#0B#),
      2063 => to_slv(opcode_type, 16#06#),
      2064 => to_slv(opcode_type, 16#09#),
      2065 => to_slv(opcode_type, 16#09#),
      2066 => to_slv(opcode_type, 16#0A#),
      2067 => to_slv(opcode_type, 16#0F#),
      2068 => to_slv(opcode_type, 16#06#),
      2069 => to_slv(opcode_type, 16#0B#),
      2070 => to_slv(opcode_type, 16#0E#),
      2071 => to_slv(opcode_type, 16#06#),
      2072 => to_slv(opcode_type, 16#08#),
      2073 => to_slv(opcode_type, 16#0E#),
      2074 => to_slv(opcode_type, 16#47#),
      2075 => to_slv(opcode_type, 16#08#),
      2076 => to_slv(opcode_type, 16#0D#),
      2077 => to_slv(opcode_type, 16#10#),
      2078 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#06#),
      2081 => to_slv(opcode_type, 16#09#),
      2082 => to_slv(opcode_type, 16#09#),
      2083 => to_slv(opcode_type, 16#03#),
      2084 => to_slv(opcode_type, 16#C8#),
      2085 => to_slv(opcode_type, 16#09#),
      2086 => to_slv(opcode_type, 16#0E#),
      2087 => to_slv(opcode_type, 16#0C#),
      2088 => to_slv(opcode_type, 16#06#),
      2089 => to_slv(opcode_type, 16#07#),
      2090 => to_slv(opcode_type, 16#11#),
      2091 => to_slv(opcode_type, 16#0C#),
      2092 => to_slv(opcode_type, 16#09#),
      2093 => to_slv(opcode_type, 16#0B#),
      2094 => to_slv(opcode_type, 16#10#),
      2095 => to_slv(opcode_type, 16#06#),
      2096 => to_slv(opcode_type, 16#07#),
      2097 => to_slv(opcode_type, 16#07#),
      2098 => to_slv(opcode_type, 16#0B#),
      2099 => to_slv(opcode_type, 16#0E#),
      2100 => to_slv(opcode_type, 16#08#),
      2101 => to_slv(opcode_type, 16#12#),
      2102 => to_slv(opcode_type, 16#23#),
      2103 => to_slv(opcode_type, 16#08#),
      2104 => to_slv(opcode_type, 16#08#),
      2105 => to_slv(opcode_type, 16#0C#),
      2106 => to_slv(opcode_type, 16#0F#),
      2107 => to_slv(opcode_type, 16#07#),
      2108 => to_slv(opcode_type, 16#11#),
      2109 => to_slv(opcode_type, 16#0E#),
      2110 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#08#),
      2113 => to_slv(opcode_type, 16#09#),
      2114 => to_slv(opcode_type, 16#06#),
      2115 => to_slv(opcode_type, 16#03#),
      2116 => to_slv(opcode_type, 16#0C#),
      2117 => to_slv(opcode_type, 16#08#),
      2118 => to_slv(opcode_type, 16#0C#),
      2119 => to_slv(opcode_type, 16#0C#),
      2120 => to_slv(opcode_type, 16#07#),
      2121 => to_slv(opcode_type, 16#07#),
      2122 => to_slv(opcode_type, 16#0B#),
      2123 => to_slv(opcode_type, 16#CE#),
      2124 => to_slv(opcode_type, 16#08#),
      2125 => to_slv(opcode_type, 16#0F#),
      2126 => to_slv(opcode_type, 16#11#),
      2127 => to_slv(opcode_type, 16#08#),
      2128 => to_slv(opcode_type, 16#06#),
      2129 => to_slv(opcode_type, 16#06#),
      2130 => to_slv(opcode_type, 16#0E#),
      2131 => to_slv(opcode_type, 16#10#),
      2132 => to_slv(opcode_type, 16#09#),
      2133 => to_slv(opcode_type, 16#0A#),
      2134 => to_slv(opcode_type, 16#0E#),
      2135 => to_slv(opcode_type, 16#06#),
      2136 => to_slv(opcode_type, 16#09#),
      2137 => to_slv(opcode_type, 16#0F#),
      2138 => to_slv(opcode_type, 16#0F#),
      2139 => to_slv(opcode_type, 16#07#),
      2140 => to_slv(opcode_type, 16#DF#),
      2141 => to_slv(opcode_type, 16#10#),
      2142 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#08#),
      2145 => to_slv(opcode_type, 16#07#),
      2146 => to_slv(opcode_type, 16#06#),
      2147 => to_slv(opcode_type, 16#02#),
      2148 => to_slv(opcode_type, 16#0E#),
      2149 => to_slv(opcode_type, 16#08#),
      2150 => to_slv(opcode_type, 16#91#),
      2151 => to_slv(opcode_type, 16#0E#),
      2152 => to_slv(opcode_type, 16#09#),
      2153 => to_slv(opcode_type, 16#08#),
      2154 => to_slv(opcode_type, 16#0D#),
      2155 => to_slv(opcode_type, 16#0C#),
      2156 => to_slv(opcode_type, 16#09#),
      2157 => to_slv(opcode_type, 16#0E#),
      2158 => to_slv(opcode_type, 16#0C#),
      2159 => to_slv(opcode_type, 16#07#),
      2160 => to_slv(opcode_type, 16#08#),
      2161 => to_slv(opcode_type, 16#06#),
      2162 => to_slv(opcode_type, 16#11#),
      2163 => to_slv(opcode_type, 16#0E#),
      2164 => to_slv(opcode_type, 16#06#),
      2165 => to_slv(opcode_type, 16#57#),
      2166 => to_slv(opcode_type, 16#0E#),
      2167 => to_slv(opcode_type, 16#07#),
      2168 => to_slv(opcode_type, 16#07#),
      2169 => to_slv(opcode_type, 16#0C#),
      2170 => to_slv(opcode_type, 16#0B#),
      2171 => to_slv(opcode_type, 16#07#),
      2172 => to_slv(opcode_type, 16#0E#),
      2173 => to_slv(opcode_type, 16#0B#),
      2174 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#07#),
      2177 => to_slv(opcode_type, 16#06#),
      2178 => to_slv(opcode_type, 16#07#),
      2179 => to_slv(opcode_type, 16#06#),
      2180 => to_slv(opcode_type, 16#10#),
      2181 => to_slv(opcode_type, 16#0E#),
      2182 => to_slv(opcode_type, 16#02#),
      2183 => to_slv(opcode_type, 16#0F#),
      2184 => to_slv(opcode_type, 16#06#),
      2185 => to_slv(opcode_type, 16#08#),
      2186 => to_slv(opcode_type, 16#0A#),
      2187 => to_slv(opcode_type, 16#0F#),
      2188 => to_slv(opcode_type, 16#08#),
      2189 => to_slv(opcode_type, 16#0A#),
      2190 => to_slv(opcode_type, 16#0D#),
      2191 => to_slv(opcode_type, 16#07#),
      2192 => to_slv(opcode_type, 16#06#),
      2193 => to_slv(opcode_type, 16#09#),
      2194 => to_slv(opcode_type, 16#11#),
      2195 => to_slv(opcode_type, 16#0C#),
      2196 => to_slv(opcode_type, 16#09#),
      2197 => to_slv(opcode_type, 16#0D#),
      2198 => to_slv(opcode_type, 16#11#),
      2199 => to_slv(opcode_type, 16#08#),
      2200 => to_slv(opcode_type, 16#07#),
      2201 => to_slv(opcode_type, 16#0C#),
      2202 => to_slv(opcode_type, 16#0F#),
      2203 => to_slv(opcode_type, 16#08#),
      2204 => to_slv(opcode_type, 16#0F#),
      2205 => to_slv(opcode_type, 16#0B#),
      2206 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#09#),
      2209 => to_slv(opcode_type, 16#06#),
      2210 => to_slv(opcode_type, 16#08#),
      2211 => to_slv(opcode_type, 16#04#),
      2212 => to_slv(opcode_type, 16#0D#),
      2213 => to_slv(opcode_type, 16#07#),
      2214 => to_slv(opcode_type, 16#0F#),
      2215 => to_slv(opcode_type, 16#0A#),
      2216 => to_slv(opcode_type, 16#07#),
      2217 => to_slv(opcode_type, 16#09#),
      2218 => to_slv(opcode_type, 16#11#),
      2219 => to_slv(opcode_type, 16#11#),
      2220 => to_slv(opcode_type, 16#09#),
      2221 => to_slv(opcode_type, 16#0B#),
      2222 => to_slv(opcode_type, 16#0B#),
      2223 => to_slv(opcode_type, 16#08#),
      2224 => to_slv(opcode_type, 16#08#),
      2225 => to_slv(opcode_type, 16#09#),
      2226 => to_slv(opcode_type, 16#11#),
      2227 => to_slv(opcode_type, 16#EC#),
      2228 => to_slv(opcode_type, 16#09#),
      2229 => to_slv(opcode_type, 16#10#),
      2230 => to_slv(opcode_type, 16#0E#),
      2231 => to_slv(opcode_type, 16#07#),
      2232 => to_slv(opcode_type, 16#07#),
      2233 => to_slv(opcode_type, 16#0B#),
      2234 => to_slv(opcode_type, 16#0F#),
      2235 => to_slv(opcode_type, 16#07#),
      2236 => to_slv(opcode_type, 16#0C#),
      2237 => to_slv(opcode_type, 16#0C#),
      2238 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#09#),
      2241 => to_slv(opcode_type, 16#07#),
      2242 => to_slv(opcode_type, 16#09#),
      2243 => to_slv(opcode_type, 16#09#),
      2244 => to_slv(opcode_type, 16#0D#),
      2245 => to_slv(opcode_type, 16#0C#),
      2246 => to_slv(opcode_type, 16#04#),
      2247 => to_slv(opcode_type, 16#0A#),
      2248 => to_slv(opcode_type, 16#09#),
      2249 => to_slv(opcode_type, 16#09#),
      2250 => to_slv(opcode_type, 16#0F#),
      2251 => to_slv(opcode_type, 16#0D#),
      2252 => to_slv(opcode_type, 16#08#),
      2253 => to_slv(opcode_type, 16#0D#),
      2254 => to_slv(opcode_type, 16#0C#),
      2255 => to_slv(opcode_type, 16#07#),
      2256 => to_slv(opcode_type, 16#08#),
      2257 => to_slv(opcode_type, 16#09#),
      2258 => to_slv(opcode_type, 16#0B#),
      2259 => to_slv(opcode_type, 16#0D#),
      2260 => to_slv(opcode_type, 16#06#),
      2261 => to_slv(opcode_type, 16#B1#),
      2262 => to_slv(opcode_type, 16#0F#),
      2263 => to_slv(opcode_type, 16#07#),
      2264 => to_slv(opcode_type, 16#09#),
      2265 => to_slv(opcode_type, 16#0B#),
      2266 => to_slv(opcode_type, 16#0E#),
      2267 => to_slv(opcode_type, 16#09#),
      2268 => to_slv(opcode_type, 16#10#),
      2269 => to_slv(opcode_type, 16#0C#),
      2270 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#09#),
      2273 => to_slv(opcode_type, 16#09#),
      2274 => to_slv(opcode_type, 16#08#),
      2275 => to_slv(opcode_type, 16#05#),
      2276 => to_slv(opcode_type, 16#0C#),
      2277 => to_slv(opcode_type, 16#08#),
      2278 => to_slv(opcode_type, 16#0E#),
      2279 => to_slv(opcode_type, 16#0D#),
      2280 => to_slv(opcode_type, 16#07#),
      2281 => to_slv(opcode_type, 16#09#),
      2282 => to_slv(opcode_type, 16#0F#),
      2283 => to_slv(opcode_type, 16#0E#),
      2284 => to_slv(opcode_type, 16#09#),
      2285 => to_slv(opcode_type, 16#0D#),
      2286 => to_slv(opcode_type, 16#0B#),
      2287 => to_slv(opcode_type, 16#08#),
      2288 => to_slv(opcode_type, 16#08#),
      2289 => to_slv(opcode_type, 16#06#),
      2290 => to_slv(opcode_type, 16#10#),
      2291 => to_slv(opcode_type, 16#10#),
      2292 => to_slv(opcode_type, 16#08#),
      2293 => to_slv(opcode_type, 16#CF#),
      2294 => to_slv(opcode_type, 16#0F#),
      2295 => to_slv(opcode_type, 16#09#),
      2296 => to_slv(opcode_type, 16#06#),
      2297 => to_slv(opcode_type, 16#0A#),
      2298 => to_slv(opcode_type, 16#0D#),
      2299 => to_slv(opcode_type, 16#07#),
      2300 => to_slv(opcode_type, 16#10#),
      2301 => to_slv(opcode_type, 16#0E#),
      2302 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#09#),
      2305 => to_slv(opcode_type, 16#08#),
      2306 => to_slv(opcode_type, 16#08#),
      2307 => to_slv(opcode_type, 16#02#),
      2308 => to_slv(opcode_type, 16#10#),
      2309 => to_slv(opcode_type, 16#08#),
      2310 => to_slv(opcode_type, 16#10#),
      2311 => to_slv(opcode_type, 16#D6#),
      2312 => to_slv(opcode_type, 16#07#),
      2313 => to_slv(opcode_type, 16#08#),
      2314 => to_slv(opcode_type, 16#10#),
      2315 => to_slv(opcode_type, 16#0C#),
      2316 => to_slv(opcode_type, 16#09#),
      2317 => to_slv(opcode_type, 16#10#),
      2318 => to_slv(opcode_type, 16#0D#),
      2319 => to_slv(opcode_type, 16#07#),
      2320 => to_slv(opcode_type, 16#08#),
      2321 => to_slv(opcode_type, 16#06#),
      2322 => to_slv(opcode_type, 16#0C#),
      2323 => to_slv(opcode_type, 16#0B#),
      2324 => to_slv(opcode_type, 16#09#),
      2325 => to_slv(opcode_type, 16#0E#),
      2326 => to_slv(opcode_type, 16#11#),
      2327 => to_slv(opcode_type, 16#06#),
      2328 => to_slv(opcode_type, 16#06#),
      2329 => to_slv(opcode_type, 16#0B#),
      2330 => to_slv(opcode_type, 16#0E#),
      2331 => to_slv(opcode_type, 16#07#),
      2332 => to_slv(opcode_type, 16#EA#),
      2333 => to_slv(opcode_type, 16#11#),
      2334 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#06#),
      2337 => to_slv(opcode_type, 16#06#),
      2338 => to_slv(opcode_type, 16#09#),
      2339 => to_slv(opcode_type, 16#01#),
      2340 => to_slv(opcode_type, 16#B8#),
      2341 => to_slv(opcode_type, 16#07#),
      2342 => to_slv(opcode_type, 16#F0#),
      2343 => to_slv(opcode_type, 16#0C#),
      2344 => to_slv(opcode_type, 16#08#),
      2345 => to_slv(opcode_type, 16#06#),
      2346 => to_slv(opcode_type, 16#0D#),
      2347 => to_slv(opcode_type, 16#0F#),
      2348 => to_slv(opcode_type, 16#08#),
      2349 => to_slv(opcode_type, 16#0A#),
      2350 => to_slv(opcode_type, 16#0F#),
      2351 => to_slv(opcode_type, 16#06#),
      2352 => to_slv(opcode_type, 16#09#),
      2353 => to_slv(opcode_type, 16#08#),
      2354 => to_slv(opcode_type, 16#0F#),
      2355 => to_slv(opcode_type, 16#0D#),
      2356 => to_slv(opcode_type, 16#06#),
      2357 => to_slv(opcode_type, 16#11#),
      2358 => to_slv(opcode_type, 16#56#),
      2359 => to_slv(opcode_type, 16#09#),
      2360 => to_slv(opcode_type, 16#09#),
      2361 => to_slv(opcode_type, 16#0E#),
      2362 => to_slv(opcode_type, 16#0E#),
      2363 => to_slv(opcode_type, 16#08#),
      2364 => to_slv(opcode_type, 16#C7#),
      2365 => to_slv(opcode_type, 16#11#),
      2366 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#08#),
      2369 => to_slv(opcode_type, 16#06#),
      2370 => to_slv(opcode_type, 16#07#),
      2371 => to_slv(opcode_type, 16#08#),
      2372 => to_slv(opcode_type, 16#11#),
      2373 => to_slv(opcode_type, 16#0B#),
      2374 => to_slv(opcode_type, 16#09#),
      2375 => to_slv(opcode_type, 16#0A#),
      2376 => to_slv(opcode_type, 16#11#),
      2377 => to_slv(opcode_type, 16#06#),
      2378 => to_slv(opcode_type, 16#04#),
      2379 => to_slv(opcode_type, 16#0A#),
      2380 => to_slv(opcode_type, 16#08#),
      2381 => to_slv(opcode_type, 16#0C#),
      2382 => to_slv(opcode_type, 16#0A#),
      2383 => to_slv(opcode_type, 16#06#),
      2384 => to_slv(opcode_type, 16#07#),
      2385 => to_slv(opcode_type, 16#09#),
      2386 => to_slv(opcode_type, 16#10#),
      2387 => to_slv(opcode_type, 16#0B#),
      2388 => to_slv(opcode_type, 16#07#),
      2389 => to_slv(opcode_type, 16#0F#),
      2390 => to_slv(opcode_type, 16#11#),
      2391 => to_slv(opcode_type, 16#09#),
      2392 => to_slv(opcode_type, 16#08#),
      2393 => to_slv(opcode_type, 16#8F#),
      2394 => to_slv(opcode_type, 16#11#),
      2395 => to_slv(opcode_type, 16#09#),
      2396 => to_slv(opcode_type, 16#0B#),
      2397 => to_slv(opcode_type, 16#3A#),
      2398 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#06#),
      2401 => to_slv(opcode_type, 16#09#),
      2402 => to_slv(opcode_type, 16#08#),
      2403 => to_slv(opcode_type, 16#09#),
      2404 => to_slv(opcode_type, 16#0A#),
      2405 => to_slv(opcode_type, 16#11#),
      2406 => to_slv(opcode_type, 16#07#),
      2407 => to_slv(opcode_type, 16#0C#),
      2408 => to_slv(opcode_type, 16#10#),
      2409 => to_slv(opcode_type, 16#06#),
      2410 => to_slv(opcode_type, 16#05#),
      2411 => to_slv(opcode_type, 16#11#),
      2412 => to_slv(opcode_type, 16#09#),
      2413 => to_slv(opcode_type, 16#10#),
      2414 => to_slv(opcode_type, 16#11#),
      2415 => to_slv(opcode_type, 16#06#),
      2416 => to_slv(opcode_type, 16#08#),
      2417 => to_slv(opcode_type, 16#07#),
      2418 => to_slv(opcode_type, 16#0A#),
      2419 => to_slv(opcode_type, 16#0F#),
      2420 => to_slv(opcode_type, 16#07#),
      2421 => to_slv(opcode_type, 16#0A#),
      2422 => to_slv(opcode_type, 16#10#),
      2423 => to_slv(opcode_type, 16#07#),
      2424 => to_slv(opcode_type, 16#09#),
      2425 => to_slv(opcode_type, 16#0D#),
      2426 => to_slv(opcode_type, 16#0B#),
      2427 => to_slv(opcode_type, 16#06#),
      2428 => to_slv(opcode_type, 16#6E#),
      2429 => to_slv(opcode_type, 16#11#),
      2430 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#06#),
      2433 => to_slv(opcode_type, 16#08#),
      2434 => to_slv(opcode_type, 16#06#),
      2435 => to_slv(opcode_type, 16#05#),
      2436 => to_slv(opcode_type, 16#0E#),
      2437 => to_slv(opcode_type, 16#07#),
      2438 => to_slv(opcode_type, 16#0D#),
      2439 => to_slv(opcode_type, 16#0D#),
      2440 => to_slv(opcode_type, 16#09#),
      2441 => to_slv(opcode_type, 16#08#),
      2442 => to_slv(opcode_type, 16#0B#),
      2443 => to_slv(opcode_type, 16#F9#),
      2444 => to_slv(opcode_type, 16#07#),
      2445 => to_slv(opcode_type, 16#0F#),
      2446 => to_slv(opcode_type, 16#97#),
      2447 => to_slv(opcode_type, 16#06#),
      2448 => to_slv(opcode_type, 16#09#),
      2449 => to_slv(opcode_type, 16#09#),
      2450 => to_slv(opcode_type, 16#0C#),
      2451 => to_slv(opcode_type, 16#10#),
      2452 => to_slv(opcode_type, 16#09#),
      2453 => to_slv(opcode_type, 16#0A#),
      2454 => to_slv(opcode_type, 16#0A#),
      2455 => to_slv(opcode_type, 16#09#),
      2456 => to_slv(opcode_type, 16#08#),
      2457 => to_slv(opcode_type, 16#0A#),
      2458 => to_slv(opcode_type, 16#0D#),
      2459 => to_slv(opcode_type, 16#08#),
      2460 => to_slv(opcode_type, 16#0B#),
      2461 => to_slv(opcode_type, 16#0F#),
      2462 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#08#),
      2465 => to_slv(opcode_type, 16#09#),
      2466 => to_slv(opcode_type, 16#09#),
      2467 => to_slv(opcode_type, 16#04#),
      2468 => to_slv(opcode_type, 16#58#),
      2469 => to_slv(opcode_type, 16#06#),
      2470 => to_slv(opcode_type, 16#11#),
      2471 => to_slv(opcode_type, 16#11#),
      2472 => to_slv(opcode_type, 16#07#),
      2473 => to_slv(opcode_type, 16#08#),
      2474 => to_slv(opcode_type, 16#11#),
      2475 => to_slv(opcode_type, 16#0A#),
      2476 => to_slv(opcode_type, 16#09#),
      2477 => to_slv(opcode_type, 16#0D#),
      2478 => to_slv(opcode_type, 16#0E#),
      2479 => to_slv(opcode_type, 16#09#),
      2480 => to_slv(opcode_type, 16#09#),
      2481 => to_slv(opcode_type, 16#09#),
      2482 => to_slv(opcode_type, 16#0A#),
      2483 => to_slv(opcode_type, 16#0D#),
      2484 => to_slv(opcode_type, 16#07#),
      2485 => to_slv(opcode_type, 16#0E#),
      2486 => to_slv(opcode_type, 16#0F#),
      2487 => to_slv(opcode_type, 16#06#),
      2488 => to_slv(opcode_type, 16#07#),
      2489 => to_slv(opcode_type, 16#0C#),
      2490 => to_slv(opcode_type, 16#0F#),
      2491 => to_slv(opcode_type, 16#08#),
      2492 => to_slv(opcode_type, 16#AC#),
      2493 => to_slv(opcode_type, 16#0A#),
      2494 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#08#),
      2497 => to_slv(opcode_type, 16#09#),
      2498 => to_slv(opcode_type, 16#09#),
      2499 => to_slv(opcode_type, 16#04#),
      2500 => to_slv(opcode_type, 16#0E#),
      2501 => to_slv(opcode_type, 16#08#),
      2502 => to_slv(opcode_type, 16#0F#),
      2503 => to_slv(opcode_type, 16#0F#),
      2504 => to_slv(opcode_type, 16#07#),
      2505 => to_slv(opcode_type, 16#07#),
      2506 => to_slv(opcode_type, 16#0E#),
      2507 => to_slv(opcode_type, 16#0F#),
      2508 => to_slv(opcode_type, 16#06#),
      2509 => to_slv(opcode_type, 16#FC#),
      2510 => to_slv(opcode_type, 16#60#),
      2511 => to_slv(opcode_type, 16#06#),
      2512 => to_slv(opcode_type, 16#09#),
      2513 => to_slv(opcode_type, 16#07#),
      2514 => to_slv(opcode_type, 16#5A#),
      2515 => to_slv(opcode_type, 16#0C#),
      2516 => to_slv(opcode_type, 16#07#),
      2517 => to_slv(opcode_type, 16#11#),
      2518 => to_slv(opcode_type, 16#0A#),
      2519 => to_slv(opcode_type, 16#09#),
      2520 => to_slv(opcode_type, 16#09#),
      2521 => to_slv(opcode_type, 16#0D#),
      2522 => to_slv(opcode_type, 16#0A#),
      2523 => to_slv(opcode_type, 16#09#),
      2524 => to_slv(opcode_type, 16#0B#),
      2525 => to_slv(opcode_type, 16#0E#),
      2526 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#08#),
      2529 => to_slv(opcode_type, 16#07#),
      2530 => to_slv(opcode_type, 16#06#),
      2531 => to_slv(opcode_type, 16#07#),
      2532 => to_slv(opcode_type, 16#0D#),
      2533 => to_slv(opcode_type, 16#0A#),
      2534 => to_slv(opcode_type, 16#01#),
      2535 => to_slv(opcode_type, 16#10#),
      2536 => to_slv(opcode_type, 16#08#),
      2537 => to_slv(opcode_type, 16#08#),
      2538 => to_slv(opcode_type, 16#0A#),
      2539 => to_slv(opcode_type, 16#0C#),
      2540 => to_slv(opcode_type, 16#08#),
      2541 => to_slv(opcode_type, 16#2C#),
      2542 => to_slv(opcode_type, 16#0D#),
      2543 => to_slv(opcode_type, 16#08#),
      2544 => to_slv(opcode_type, 16#09#),
      2545 => to_slv(opcode_type, 16#08#),
      2546 => to_slv(opcode_type, 16#11#),
      2547 => to_slv(opcode_type, 16#0F#),
      2548 => to_slv(opcode_type, 16#06#),
      2549 => to_slv(opcode_type, 16#0C#),
      2550 => to_slv(opcode_type, 16#10#),
      2551 => to_slv(opcode_type, 16#07#),
      2552 => to_slv(opcode_type, 16#09#),
      2553 => to_slv(opcode_type, 16#10#),
      2554 => to_slv(opcode_type, 16#0B#),
      2555 => to_slv(opcode_type, 16#08#),
      2556 => to_slv(opcode_type, 16#0C#),
      2557 => to_slv(opcode_type, 16#0A#),
      2558 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#09#),
      2561 => to_slv(opcode_type, 16#09#),
      2562 => to_slv(opcode_type, 16#08#),
      2563 => to_slv(opcode_type, 16#03#),
      2564 => to_slv(opcode_type, 16#11#),
      2565 => to_slv(opcode_type, 16#06#),
      2566 => to_slv(opcode_type, 16#11#),
      2567 => to_slv(opcode_type, 16#0F#),
      2568 => to_slv(opcode_type, 16#07#),
      2569 => to_slv(opcode_type, 16#07#),
      2570 => to_slv(opcode_type, 16#0D#),
      2571 => to_slv(opcode_type, 16#11#),
      2572 => to_slv(opcode_type, 16#06#),
      2573 => to_slv(opcode_type, 16#0E#),
      2574 => to_slv(opcode_type, 16#11#),
      2575 => to_slv(opcode_type, 16#07#),
      2576 => to_slv(opcode_type, 16#09#),
      2577 => to_slv(opcode_type, 16#08#),
      2578 => to_slv(opcode_type, 16#0E#),
      2579 => to_slv(opcode_type, 16#0D#),
      2580 => to_slv(opcode_type, 16#07#),
      2581 => to_slv(opcode_type, 16#0B#),
      2582 => to_slv(opcode_type, 16#11#),
      2583 => to_slv(opcode_type, 16#09#),
      2584 => to_slv(opcode_type, 16#09#),
      2585 => to_slv(opcode_type, 16#0F#),
      2586 => to_slv(opcode_type, 16#0C#),
      2587 => to_slv(opcode_type, 16#07#),
      2588 => to_slv(opcode_type, 16#11#),
      2589 => to_slv(opcode_type, 16#0A#),
      2590 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#09#),
      2593 => to_slv(opcode_type, 16#07#),
      2594 => to_slv(opcode_type, 16#06#),
      2595 => to_slv(opcode_type, 16#01#),
      2596 => to_slv(opcode_type, 16#10#),
      2597 => to_slv(opcode_type, 16#06#),
      2598 => to_slv(opcode_type, 16#0B#),
      2599 => to_slv(opcode_type, 16#10#),
      2600 => to_slv(opcode_type, 16#08#),
      2601 => to_slv(opcode_type, 16#08#),
      2602 => to_slv(opcode_type, 16#0E#),
      2603 => to_slv(opcode_type, 16#0E#),
      2604 => to_slv(opcode_type, 16#09#),
      2605 => to_slv(opcode_type, 16#11#),
      2606 => to_slv(opcode_type, 16#0D#),
      2607 => to_slv(opcode_type, 16#08#),
      2608 => to_slv(opcode_type, 16#08#),
      2609 => to_slv(opcode_type, 16#06#),
      2610 => to_slv(opcode_type, 16#0E#),
      2611 => to_slv(opcode_type, 16#0C#),
      2612 => to_slv(opcode_type, 16#07#),
      2613 => to_slv(opcode_type, 16#0A#),
      2614 => to_slv(opcode_type, 16#0D#),
      2615 => to_slv(opcode_type, 16#06#),
      2616 => to_slv(opcode_type, 16#06#),
      2617 => to_slv(opcode_type, 16#0F#),
      2618 => to_slv(opcode_type, 16#0E#),
      2619 => to_slv(opcode_type, 16#09#),
      2620 => to_slv(opcode_type, 16#0B#),
      2621 => to_slv(opcode_type, 16#0C#),
      2622 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#09#),
      2625 => to_slv(opcode_type, 16#07#),
      2626 => to_slv(opcode_type, 16#07#),
      2627 => to_slv(opcode_type, 16#06#),
      2628 => to_slv(opcode_type, 16#11#),
      2629 => to_slv(opcode_type, 16#0A#),
      2630 => to_slv(opcode_type, 16#07#),
      2631 => to_slv(opcode_type, 16#11#),
      2632 => to_slv(opcode_type, 16#0E#),
      2633 => to_slv(opcode_type, 16#09#),
      2634 => to_slv(opcode_type, 16#07#),
      2635 => to_slv(opcode_type, 16#0A#),
      2636 => to_slv(opcode_type, 16#0C#),
      2637 => to_slv(opcode_type, 16#02#),
      2638 => to_slv(opcode_type, 16#0E#),
      2639 => to_slv(opcode_type, 16#06#),
      2640 => to_slv(opcode_type, 16#09#),
      2641 => to_slv(opcode_type, 16#08#),
      2642 => to_slv(opcode_type, 16#0D#),
      2643 => to_slv(opcode_type, 16#0C#),
      2644 => to_slv(opcode_type, 16#08#),
      2645 => to_slv(opcode_type, 16#11#),
      2646 => to_slv(opcode_type, 16#D6#),
      2647 => to_slv(opcode_type, 16#09#),
      2648 => to_slv(opcode_type, 16#06#),
      2649 => to_slv(opcode_type, 16#C5#),
      2650 => to_slv(opcode_type, 16#0F#),
      2651 => to_slv(opcode_type, 16#06#),
      2652 => to_slv(opcode_type, 16#10#),
      2653 => to_slv(opcode_type, 16#11#),
      2654 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#06#),
      2657 => to_slv(opcode_type, 16#06#),
      2658 => to_slv(opcode_type, 16#07#),
      2659 => to_slv(opcode_type, 16#01#),
      2660 => to_slv(opcode_type, 16#0C#),
      2661 => to_slv(opcode_type, 16#07#),
      2662 => to_slv(opcode_type, 16#0E#),
      2663 => to_slv(opcode_type, 16#0F#),
      2664 => to_slv(opcode_type, 16#07#),
      2665 => to_slv(opcode_type, 16#07#),
      2666 => to_slv(opcode_type, 16#11#),
      2667 => to_slv(opcode_type, 16#0D#),
      2668 => to_slv(opcode_type, 16#09#),
      2669 => to_slv(opcode_type, 16#0B#),
      2670 => to_slv(opcode_type, 16#0F#),
      2671 => to_slv(opcode_type, 16#07#),
      2672 => to_slv(opcode_type, 16#09#),
      2673 => to_slv(opcode_type, 16#07#),
      2674 => to_slv(opcode_type, 16#0D#),
      2675 => to_slv(opcode_type, 16#0B#),
      2676 => to_slv(opcode_type, 16#09#),
      2677 => to_slv(opcode_type, 16#0A#),
      2678 => to_slv(opcode_type, 16#11#),
      2679 => to_slv(opcode_type, 16#07#),
      2680 => to_slv(opcode_type, 16#08#),
      2681 => to_slv(opcode_type, 16#AD#),
      2682 => to_slv(opcode_type, 16#10#),
      2683 => to_slv(opcode_type, 16#07#),
      2684 => to_slv(opcode_type, 16#0D#),
      2685 => to_slv(opcode_type, 16#D2#),
      2686 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#09#),
      2689 => to_slv(opcode_type, 16#06#),
      2690 => to_slv(opcode_type, 16#08#),
      2691 => to_slv(opcode_type, 16#07#),
      2692 => to_slv(opcode_type, 16#0F#),
      2693 => to_slv(opcode_type, 16#AB#),
      2694 => to_slv(opcode_type, 16#07#),
      2695 => to_slv(opcode_type, 16#11#),
      2696 => to_slv(opcode_type, 16#11#),
      2697 => to_slv(opcode_type, 16#08#),
      2698 => to_slv(opcode_type, 16#03#),
      2699 => to_slv(opcode_type, 16#0E#),
      2700 => to_slv(opcode_type, 16#08#),
      2701 => to_slv(opcode_type, 16#10#),
      2702 => to_slv(opcode_type, 16#11#),
      2703 => to_slv(opcode_type, 16#07#),
      2704 => to_slv(opcode_type, 16#06#),
      2705 => to_slv(opcode_type, 16#09#),
      2706 => to_slv(opcode_type, 16#D6#),
      2707 => to_slv(opcode_type, 16#11#),
      2708 => to_slv(opcode_type, 16#08#),
      2709 => to_slv(opcode_type, 16#11#),
      2710 => to_slv(opcode_type, 16#11#),
      2711 => to_slv(opcode_type, 16#07#),
      2712 => to_slv(opcode_type, 16#09#),
      2713 => to_slv(opcode_type, 16#0D#),
      2714 => to_slv(opcode_type, 16#DD#),
      2715 => to_slv(opcode_type, 16#08#),
      2716 => to_slv(opcode_type, 16#11#),
      2717 => to_slv(opcode_type, 16#11#),
      2718 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#08#),
      2721 => to_slv(opcode_type, 16#07#),
      2722 => to_slv(opcode_type, 16#08#),
      2723 => to_slv(opcode_type, 16#06#),
      2724 => to_slv(opcode_type, 16#0A#),
      2725 => to_slv(opcode_type, 16#2B#),
      2726 => to_slv(opcode_type, 16#07#),
      2727 => to_slv(opcode_type, 16#11#),
      2728 => to_slv(opcode_type, 16#A7#),
      2729 => to_slv(opcode_type, 16#07#),
      2730 => to_slv(opcode_type, 16#09#),
      2731 => to_slv(opcode_type, 16#90#),
      2732 => to_slv(opcode_type, 16#10#),
      2733 => to_slv(opcode_type, 16#08#),
      2734 => to_slv(opcode_type, 16#0F#),
      2735 => to_slv(opcode_type, 16#0B#),
      2736 => to_slv(opcode_type, 16#06#),
      2737 => to_slv(opcode_type, 16#08#),
      2738 => to_slv(opcode_type, 16#04#),
      2739 => to_slv(opcode_type, 16#0E#),
      2740 => to_slv(opcode_type, 16#06#),
      2741 => to_slv(opcode_type, 16#11#),
      2742 => to_slv(opcode_type, 16#0C#),
      2743 => to_slv(opcode_type, 16#09#),
      2744 => to_slv(opcode_type, 16#06#),
      2745 => to_slv(opcode_type, 16#0B#),
      2746 => to_slv(opcode_type, 16#0E#),
      2747 => to_slv(opcode_type, 16#07#),
      2748 => to_slv(opcode_type, 16#11#),
      2749 => to_slv(opcode_type, 16#0F#),
      2750 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#08#),
      2753 => to_slv(opcode_type, 16#09#),
      2754 => to_slv(opcode_type, 16#09#),
      2755 => to_slv(opcode_type, 16#03#),
      2756 => to_slv(opcode_type, 16#10#),
      2757 => to_slv(opcode_type, 16#06#),
      2758 => to_slv(opcode_type, 16#0E#),
      2759 => to_slv(opcode_type, 16#0E#),
      2760 => to_slv(opcode_type, 16#06#),
      2761 => to_slv(opcode_type, 16#07#),
      2762 => to_slv(opcode_type, 16#0D#),
      2763 => to_slv(opcode_type, 16#0B#),
      2764 => to_slv(opcode_type, 16#06#),
      2765 => to_slv(opcode_type, 16#0C#),
      2766 => to_slv(opcode_type, 16#10#),
      2767 => to_slv(opcode_type, 16#07#),
      2768 => to_slv(opcode_type, 16#07#),
      2769 => to_slv(opcode_type, 16#09#),
      2770 => to_slv(opcode_type, 16#11#),
      2771 => to_slv(opcode_type, 16#0C#),
      2772 => to_slv(opcode_type, 16#06#),
      2773 => to_slv(opcode_type, 16#11#),
      2774 => to_slv(opcode_type, 16#11#),
      2775 => to_slv(opcode_type, 16#07#),
      2776 => to_slv(opcode_type, 16#06#),
      2777 => to_slv(opcode_type, 16#0B#),
      2778 => to_slv(opcode_type, 16#0B#),
      2779 => to_slv(opcode_type, 16#08#),
      2780 => to_slv(opcode_type, 16#0A#),
      2781 => to_slv(opcode_type, 16#0B#),
      2782 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#09#),
      2785 => to_slv(opcode_type, 16#07#),
      2786 => to_slv(opcode_type, 16#07#),
      2787 => to_slv(opcode_type, 16#04#),
      2788 => to_slv(opcode_type, 16#0B#),
      2789 => to_slv(opcode_type, 16#06#),
      2790 => to_slv(opcode_type, 16#11#),
      2791 => to_slv(opcode_type, 16#10#),
      2792 => to_slv(opcode_type, 16#07#),
      2793 => to_slv(opcode_type, 16#08#),
      2794 => to_slv(opcode_type, 16#10#),
      2795 => to_slv(opcode_type, 16#0A#),
      2796 => to_slv(opcode_type, 16#07#),
      2797 => to_slv(opcode_type, 16#0F#),
      2798 => to_slv(opcode_type, 16#0E#),
      2799 => to_slv(opcode_type, 16#06#),
      2800 => to_slv(opcode_type, 16#09#),
      2801 => to_slv(opcode_type, 16#09#),
      2802 => to_slv(opcode_type, 16#F7#),
      2803 => to_slv(opcode_type, 16#11#),
      2804 => to_slv(opcode_type, 16#06#),
      2805 => to_slv(opcode_type, 16#0F#),
      2806 => to_slv(opcode_type, 16#0B#),
      2807 => to_slv(opcode_type, 16#08#),
      2808 => to_slv(opcode_type, 16#08#),
      2809 => to_slv(opcode_type, 16#10#),
      2810 => to_slv(opcode_type, 16#0D#),
      2811 => to_slv(opcode_type, 16#08#),
      2812 => to_slv(opcode_type, 16#0F#),
      2813 => to_slv(opcode_type, 16#0A#),
      2814 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#06#),
      2817 => to_slv(opcode_type, 16#09#),
      2818 => to_slv(opcode_type, 16#06#),
      2819 => to_slv(opcode_type, 16#05#),
      2820 => to_slv(opcode_type, 16#0E#),
      2821 => to_slv(opcode_type, 16#08#),
      2822 => to_slv(opcode_type, 16#0B#),
      2823 => to_slv(opcode_type, 16#0B#),
      2824 => to_slv(opcode_type, 16#08#),
      2825 => to_slv(opcode_type, 16#07#),
      2826 => to_slv(opcode_type, 16#0A#),
      2827 => to_slv(opcode_type, 16#0C#),
      2828 => to_slv(opcode_type, 16#09#),
      2829 => to_slv(opcode_type, 16#0E#),
      2830 => to_slv(opcode_type, 16#0F#),
      2831 => to_slv(opcode_type, 16#08#),
      2832 => to_slv(opcode_type, 16#07#),
      2833 => to_slv(opcode_type, 16#06#),
      2834 => to_slv(opcode_type, 16#0B#),
      2835 => to_slv(opcode_type, 16#0A#),
      2836 => to_slv(opcode_type, 16#07#),
      2837 => to_slv(opcode_type, 16#0F#),
      2838 => to_slv(opcode_type, 16#0B#),
      2839 => to_slv(opcode_type, 16#07#),
      2840 => to_slv(opcode_type, 16#06#),
      2841 => to_slv(opcode_type, 16#10#),
      2842 => to_slv(opcode_type, 16#5C#),
      2843 => to_slv(opcode_type, 16#09#),
      2844 => to_slv(opcode_type, 16#0D#),
      2845 => to_slv(opcode_type, 16#0C#),
      2846 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#07#),
      2849 => to_slv(opcode_type, 16#09#),
      2850 => to_slv(opcode_type, 16#08#),
      2851 => to_slv(opcode_type, 16#01#),
      2852 => to_slv(opcode_type, 16#0E#),
      2853 => to_slv(opcode_type, 16#09#),
      2854 => to_slv(opcode_type, 16#10#),
      2855 => to_slv(opcode_type, 16#0E#),
      2856 => to_slv(opcode_type, 16#09#),
      2857 => to_slv(opcode_type, 16#07#),
      2858 => to_slv(opcode_type, 16#0A#),
      2859 => to_slv(opcode_type, 16#0A#),
      2860 => to_slv(opcode_type, 16#06#),
      2861 => to_slv(opcode_type, 16#0F#),
      2862 => to_slv(opcode_type, 16#0F#),
      2863 => to_slv(opcode_type, 16#06#),
      2864 => to_slv(opcode_type, 16#06#),
      2865 => to_slv(opcode_type, 16#09#),
      2866 => to_slv(opcode_type, 16#0E#),
      2867 => to_slv(opcode_type, 16#10#),
      2868 => to_slv(opcode_type, 16#06#),
      2869 => to_slv(opcode_type, 16#0F#),
      2870 => to_slv(opcode_type, 16#0C#),
      2871 => to_slv(opcode_type, 16#07#),
      2872 => to_slv(opcode_type, 16#07#),
      2873 => to_slv(opcode_type, 16#0B#),
      2874 => to_slv(opcode_type, 16#11#),
      2875 => to_slv(opcode_type, 16#09#),
      2876 => to_slv(opcode_type, 16#0C#),
      2877 => to_slv(opcode_type, 16#11#),
      2878 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#09#),
      2881 => to_slv(opcode_type, 16#07#),
      2882 => to_slv(opcode_type, 16#06#),
      2883 => to_slv(opcode_type, 16#08#),
      2884 => to_slv(opcode_type, 16#0A#),
      2885 => to_slv(opcode_type, 16#CB#),
      2886 => to_slv(opcode_type, 16#08#),
      2887 => to_slv(opcode_type, 16#0E#),
      2888 => to_slv(opcode_type, 16#0F#),
      2889 => to_slv(opcode_type, 16#06#),
      2890 => to_slv(opcode_type, 16#07#),
      2891 => to_slv(opcode_type, 16#11#),
      2892 => to_slv(opcode_type, 16#0A#),
      2893 => to_slv(opcode_type, 16#08#),
      2894 => to_slv(opcode_type, 16#0A#),
      2895 => to_slv(opcode_type, 16#0F#),
      2896 => to_slv(opcode_type, 16#08#),
      2897 => to_slv(opcode_type, 16#06#),
      2898 => to_slv(opcode_type, 16#02#),
      2899 => to_slv(opcode_type, 16#0C#),
      2900 => to_slv(opcode_type, 16#09#),
      2901 => to_slv(opcode_type, 16#10#),
      2902 => to_slv(opcode_type, 16#BB#),
      2903 => to_slv(opcode_type, 16#08#),
      2904 => to_slv(opcode_type, 16#08#),
      2905 => to_slv(opcode_type, 16#8B#),
      2906 => to_slv(opcode_type, 16#0D#),
      2907 => to_slv(opcode_type, 16#07#),
      2908 => to_slv(opcode_type, 16#11#),
      2909 => to_slv(opcode_type, 16#0E#),
      2910 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#09#),
      2913 => to_slv(opcode_type, 16#08#),
      2914 => to_slv(opcode_type, 16#07#),
      2915 => to_slv(opcode_type, 16#09#),
      2916 => to_slv(opcode_type, 16#11#),
      2917 => to_slv(opcode_type, 16#0B#),
      2918 => to_slv(opcode_type, 16#06#),
      2919 => to_slv(opcode_type, 16#0C#),
      2920 => to_slv(opcode_type, 16#0A#),
      2921 => to_slv(opcode_type, 16#07#),
      2922 => to_slv(opcode_type, 16#06#),
      2923 => to_slv(opcode_type, 16#0E#),
      2924 => to_slv(opcode_type, 16#0C#),
      2925 => to_slv(opcode_type, 16#07#),
      2926 => to_slv(opcode_type, 16#0B#),
      2927 => to_slv(opcode_type, 16#0C#),
      2928 => to_slv(opcode_type, 16#07#),
      2929 => to_slv(opcode_type, 16#06#),
      2930 => to_slv(opcode_type, 16#08#),
      2931 => to_slv(opcode_type, 16#0A#),
      2932 => to_slv(opcode_type, 16#0A#),
      2933 => to_slv(opcode_type, 16#05#),
      2934 => to_slv(opcode_type, 16#0A#),
      2935 => to_slv(opcode_type, 16#06#),
      2936 => to_slv(opcode_type, 16#09#),
      2937 => to_slv(opcode_type, 16#0D#),
      2938 => to_slv(opcode_type, 16#0E#),
      2939 => to_slv(opcode_type, 16#08#),
      2940 => to_slv(opcode_type, 16#0A#),
      2941 => to_slv(opcode_type, 16#11#),
      2942 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#08#),
      2945 => to_slv(opcode_type, 16#06#),
      2946 => to_slv(opcode_type, 16#07#),
      2947 => to_slv(opcode_type, 16#08#),
      2948 => to_slv(opcode_type, 16#0A#),
      2949 => to_slv(opcode_type, 16#0A#),
      2950 => to_slv(opcode_type, 16#01#),
      2951 => to_slv(opcode_type, 16#0D#),
      2952 => to_slv(opcode_type, 16#07#),
      2953 => to_slv(opcode_type, 16#07#),
      2954 => to_slv(opcode_type, 16#0D#),
      2955 => to_slv(opcode_type, 16#0D#),
      2956 => to_slv(opcode_type, 16#06#),
      2957 => to_slv(opcode_type, 16#0A#),
      2958 => to_slv(opcode_type, 16#10#),
      2959 => to_slv(opcode_type, 16#07#),
      2960 => to_slv(opcode_type, 16#09#),
      2961 => to_slv(opcode_type, 16#07#),
      2962 => to_slv(opcode_type, 16#52#),
      2963 => to_slv(opcode_type, 16#0D#),
      2964 => to_slv(opcode_type, 16#08#),
      2965 => to_slv(opcode_type, 16#0C#),
      2966 => to_slv(opcode_type, 16#6D#),
      2967 => to_slv(opcode_type, 16#06#),
      2968 => to_slv(opcode_type, 16#08#),
      2969 => to_slv(opcode_type, 16#11#),
      2970 => to_slv(opcode_type, 16#0F#),
      2971 => to_slv(opcode_type, 16#08#),
      2972 => to_slv(opcode_type, 16#0E#),
      2973 => to_slv(opcode_type, 16#10#),
      2974 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#07#),
      2977 => to_slv(opcode_type, 16#07#),
      2978 => to_slv(opcode_type, 16#07#),
      2979 => to_slv(opcode_type, 16#05#),
      2980 => to_slv(opcode_type, 16#0D#),
      2981 => to_slv(opcode_type, 16#09#),
      2982 => to_slv(opcode_type, 16#10#),
      2983 => to_slv(opcode_type, 16#11#),
      2984 => to_slv(opcode_type, 16#07#),
      2985 => to_slv(opcode_type, 16#08#),
      2986 => to_slv(opcode_type, 16#0F#),
      2987 => to_slv(opcode_type, 16#D4#),
      2988 => to_slv(opcode_type, 16#06#),
      2989 => to_slv(opcode_type, 16#11#),
      2990 => to_slv(opcode_type, 16#11#),
      2991 => to_slv(opcode_type, 16#09#),
      2992 => to_slv(opcode_type, 16#06#),
      2993 => to_slv(opcode_type, 16#09#),
      2994 => to_slv(opcode_type, 16#0B#),
      2995 => to_slv(opcode_type, 16#0B#),
      2996 => to_slv(opcode_type, 16#08#),
      2997 => to_slv(opcode_type, 16#10#),
      2998 => to_slv(opcode_type, 16#DF#),
      2999 => to_slv(opcode_type, 16#08#),
      3000 => to_slv(opcode_type, 16#06#),
      3001 => to_slv(opcode_type, 16#0A#),
      3002 => to_slv(opcode_type, 16#11#),
      3003 => to_slv(opcode_type, 16#06#),
      3004 => to_slv(opcode_type, 16#11#),
      3005 => to_slv(opcode_type, 16#B1#),
      3006 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#08#),
      3009 => to_slv(opcode_type, 16#07#),
      3010 => to_slv(opcode_type, 16#06#),
      3011 => to_slv(opcode_type, 16#04#),
      3012 => to_slv(opcode_type, 16#11#),
      3013 => to_slv(opcode_type, 16#08#),
      3014 => to_slv(opcode_type, 16#10#),
      3015 => to_slv(opcode_type, 16#0B#),
      3016 => to_slv(opcode_type, 16#09#),
      3017 => to_slv(opcode_type, 16#07#),
      3018 => to_slv(opcode_type, 16#10#),
      3019 => to_slv(opcode_type, 16#10#),
      3020 => to_slv(opcode_type, 16#08#),
      3021 => to_slv(opcode_type, 16#0F#),
      3022 => to_slv(opcode_type, 16#0E#),
      3023 => to_slv(opcode_type, 16#08#),
      3024 => to_slv(opcode_type, 16#06#),
      3025 => to_slv(opcode_type, 16#07#),
      3026 => to_slv(opcode_type, 16#0B#),
      3027 => to_slv(opcode_type, 16#0D#),
      3028 => to_slv(opcode_type, 16#08#),
      3029 => to_slv(opcode_type, 16#0A#),
      3030 => to_slv(opcode_type, 16#0F#),
      3031 => to_slv(opcode_type, 16#06#),
      3032 => to_slv(opcode_type, 16#09#),
      3033 => to_slv(opcode_type, 16#0F#),
      3034 => to_slv(opcode_type, 16#0E#),
      3035 => to_slv(opcode_type, 16#08#),
      3036 => to_slv(opcode_type, 16#0D#),
      3037 => to_slv(opcode_type, 16#0E#),
      3038 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#09#),
      3041 => to_slv(opcode_type, 16#08#),
      3042 => to_slv(opcode_type, 16#08#),
      3043 => to_slv(opcode_type, 16#09#),
      3044 => to_slv(opcode_type, 16#0B#),
      3045 => to_slv(opcode_type, 16#0B#),
      3046 => to_slv(opcode_type, 16#02#),
      3047 => to_slv(opcode_type, 16#0F#),
      3048 => to_slv(opcode_type, 16#07#),
      3049 => to_slv(opcode_type, 16#09#),
      3050 => to_slv(opcode_type, 16#EC#),
      3051 => to_slv(opcode_type, 16#11#),
      3052 => to_slv(opcode_type, 16#07#),
      3053 => to_slv(opcode_type, 16#D7#),
      3054 => to_slv(opcode_type, 16#48#),
      3055 => to_slv(opcode_type, 16#09#),
      3056 => to_slv(opcode_type, 16#07#),
      3057 => to_slv(opcode_type, 16#09#),
      3058 => to_slv(opcode_type, 16#0E#),
      3059 => to_slv(opcode_type, 16#CF#),
      3060 => to_slv(opcode_type, 16#08#),
      3061 => to_slv(opcode_type, 16#0C#),
      3062 => to_slv(opcode_type, 16#0A#),
      3063 => to_slv(opcode_type, 16#07#),
      3064 => to_slv(opcode_type, 16#06#),
      3065 => to_slv(opcode_type, 16#0F#),
      3066 => to_slv(opcode_type, 16#0B#),
      3067 => to_slv(opcode_type, 16#07#),
      3068 => to_slv(opcode_type, 16#0A#),
      3069 => to_slv(opcode_type, 16#1F#),
      3070 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#08#),
      3073 => to_slv(opcode_type, 16#06#),
      3074 => to_slv(opcode_type, 16#06#),
      3075 => to_slv(opcode_type, 16#05#),
      3076 => to_slv(opcode_type, 16#0A#),
      3077 => to_slv(opcode_type, 16#09#),
      3078 => to_slv(opcode_type, 16#11#),
      3079 => to_slv(opcode_type, 16#0E#),
      3080 => to_slv(opcode_type, 16#06#),
      3081 => to_slv(opcode_type, 16#08#),
      3082 => to_slv(opcode_type, 16#6B#),
      3083 => to_slv(opcode_type, 16#0A#),
      3084 => to_slv(opcode_type, 16#09#),
      3085 => to_slv(opcode_type, 16#0E#),
      3086 => to_slv(opcode_type, 16#0D#),
      3087 => to_slv(opcode_type, 16#09#),
      3088 => to_slv(opcode_type, 16#09#),
      3089 => to_slv(opcode_type, 16#07#),
      3090 => to_slv(opcode_type, 16#0A#),
      3091 => to_slv(opcode_type, 16#0B#),
      3092 => to_slv(opcode_type, 16#06#),
      3093 => to_slv(opcode_type, 16#0A#),
      3094 => to_slv(opcode_type, 16#0E#),
      3095 => to_slv(opcode_type, 16#07#),
      3096 => to_slv(opcode_type, 16#09#),
      3097 => to_slv(opcode_type, 16#17#),
      3098 => to_slv(opcode_type, 16#0F#),
      3099 => to_slv(opcode_type, 16#07#),
      3100 => to_slv(opcode_type, 16#0A#),
      3101 => to_slv(opcode_type, 16#0B#),
      3102 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#08#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#06#),
      3107 => to_slv(opcode_type, 16#01#),
      3108 => to_slv(opcode_type, 16#6B#),
      3109 => to_slv(opcode_type, 16#09#),
      3110 => to_slv(opcode_type, 16#4F#),
      3111 => to_slv(opcode_type, 16#0F#),
      3112 => to_slv(opcode_type, 16#08#),
      3113 => to_slv(opcode_type, 16#08#),
      3114 => to_slv(opcode_type, 16#10#),
      3115 => to_slv(opcode_type, 16#0B#),
      3116 => to_slv(opcode_type, 16#07#),
      3117 => to_slv(opcode_type, 16#0F#),
      3118 => to_slv(opcode_type, 16#11#),
      3119 => to_slv(opcode_type, 16#06#),
      3120 => to_slv(opcode_type, 16#08#),
      3121 => to_slv(opcode_type, 16#06#),
      3122 => to_slv(opcode_type, 16#B6#),
      3123 => to_slv(opcode_type, 16#0F#),
      3124 => to_slv(opcode_type, 16#08#),
      3125 => to_slv(opcode_type, 16#0D#),
      3126 => to_slv(opcode_type, 16#0A#),
      3127 => to_slv(opcode_type, 16#09#),
      3128 => to_slv(opcode_type, 16#06#),
      3129 => to_slv(opcode_type, 16#0F#),
      3130 => to_slv(opcode_type, 16#0A#),
      3131 => to_slv(opcode_type, 16#09#),
      3132 => to_slv(opcode_type, 16#0C#),
      3133 => to_slv(opcode_type, 16#0E#),
      3134 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#09#),
      3137 => to_slv(opcode_type, 16#06#),
      3138 => to_slv(opcode_type, 16#07#),
      3139 => to_slv(opcode_type, 16#06#),
      3140 => to_slv(opcode_type, 16#10#),
      3141 => to_slv(opcode_type, 16#0A#),
      3142 => to_slv(opcode_type, 16#03#),
      3143 => to_slv(opcode_type, 16#0C#),
      3144 => to_slv(opcode_type, 16#07#),
      3145 => to_slv(opcode_type, 16#07#),
      3146 => to_slv(opcode_type, 16#0A#),
      3147 => to_slv(opcode_type, 16#0A#),
      3148 => to_slv(opcode_type, 16#07#),
      3149 => to_slv(opcode_type, 16#0E#),
      3150 => to_slv(opcode_type, 16#0B#),
      3151 => to_slv(opcode_type, 16#08#),
      3152 => to_slv(opcode_type, 16#09#),
      3153 => to_slv(opcode_type, 16#07#),
      3154 => to_slv(opcode_type, 16#0F#),
      3155 => to_slv(opcode_type, 16#0D#),
      3156 => to_slv(opcode_type, 16#08#),
      3157 => to_slv(opcode_type, 16#0E#),
      3158 => to_slv(opcode_type, 16#0D#),
      3159 => to_slv(opcode_type, 16#08#),
      3160 => to_slv(opcode_type, 16#07#),
      3161 => to_slv(opcode_type, 16#0C#),
      3162 => to_slv(opcode_type, 16#0E#),
      3163 => to_slv(opcode_type, 16#06#),
      3164 => to_slv(opcode_type, 16#0D#),
      3165 => to_slv(opcode_type, 16#0F#),
      3166 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#06#),
      3169 => to_slv(opcode_type, 16#06#),
      3170 => to_slv(opcode_type, 16#09#),
      3171 => to_slv(opcode_type, 16#07#),
      3172 => to_slv(opcode_type, 16#10#),
      3173 => to_slv(opcode_type, 16#0F#),
      3174 => to_slv(opcode_type, 16#04#),
      3175 => to_slv(opcode_type, 16#0B#),
      3176 => to_slv(opcode_type, 16#09#),
      3177 => to_slv(opcode_type, 16#09#),
      3178 => to_slv(opcode_type, 16#0D#),
      3179 => to_slv(opcode_type, 16#10#),
      3180 => to_slv(opcode_type, 16#08#),
      3181 => to_slv(opcode_type, 16#0B#),
      3182 => to_slv(opcode_type, 16#0F#),
      3183 => to_slv(opcode_type, 16#09#),
      3184 => to_slv(opcode_type, 16#09#),
      3185 => to_slv(opcode_type, 16#07#),
      3186 => to_slv(opcode_type, 16#0D#),
      3187 => to_slv(opcode_type, 16#0B#),
      3188 => to_slv(opcode_type, 16#08#),
      3189 => to_slv(opcode_type, 16#0A#),
      3190 => to_slv(opcode_type, 16#10#),
      3191 => to_slv(opcode_type, 16#09#),
      3192 => to_slv(opcode_type, 16#06#),
      3193 => to_slv(opcode_type, 16#0B#),
      3194 => to_slv(opcode_type, 16#0A#),
      3195 => to_slv(opcode_type, 16#07#),
      3196 => to_slv(opcode_type, 16#0E#),
      3197 => to_slv(opcode_type, 16#0D#),
      3198 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#06#),
      3201 => to_slv(opcode_type, 16#06#),
      3202 => to_slv(opcode_type, 16#08#),
      3203 => to_slv(opcode_type, 16#09#),
      3204 => to_slv(opcode_type, 16#0B#),
      3205 => to_slv(opcode_type, 16#0D#),
      3206 => to_slv(opcode_type, 16#03#),
      3207 => to_slv(opcode_type, 16#0A#),
      3208 => to_slv(opcode_type, 16#06#),
      3209 => to_slv(opcode_type, 16#06#),
      3210 => to_slv(opcode_type, 16#10#),
      3211 => to_slv(opcode_type, 16#0F#),
      3212 => to_slv(opcode_type, 16#09#),
      3213 => to_slv(opcode_type, 16#0A#),
      3214 => to_slv(opcode_type, 16#0A#),
      3215 => to_slv(opcode_type, 16#08#),
      3216 => to_slv(opcode_type, 16#06#),
      3217 => to_slv(opcode_type, 16#09#),
      3218 => to_slv(opcode_type, 16#11#),
      3219 => to_slv(opcode_type, 16#0C#),
      3220 => to_slv(opcode_type, 16#08#),
      3221 => to_slv(opcode_type, 16#0A#),
      3222 => to_slv(opcode_type, 16#0E#),
      3223 => to_slv(opcode_type, 16#08#),
      3224 => to_slv(opcode_type, 16#09#),
      3225 => to_slv(opcode_type, 16#3E#),
      3226 => to_slv(opcode_type, 16#0D#),
      3227 => to_slv(opcode_type, 16#09#),
      3228 => to_slv(opcode_type, 16#4A#),
      3229 => to_slv(opcode_type, 16#10#),
      3230 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#06#),
      3233 => to_slv(opcode_type, 16#09#),
      3234 => to_slv(opcode_type, 16#06#),
      3235 => to_slv(opcode_type, 16#06#),
      3236 => to_slv(opcode_type, 16#0F#),
      3237 => to_slv(opcode_type, 16#0C#),
      3238 => to_slv(opcode_type, 16#07#),
      3239 => to_slv(opcode_type, 16#0E#),
      3240 => to_slv(opcode_type, 16#0F#),
      3241 => to_slv(opcode_type, 16#06#),
      3242 => to_slv(opcode_type, 16#01#),
      3243 => to_slv(opcode_type, 16#0E#),
      3244 => to_slv(opcode_type, 16#06#),
      3245 => to_slv(opcode_type, 16#11#),
      3246 => to_slv(opcode_type, 16#0C#),
      3247 => to_slv(opcode_type, 16#06#),
      3248 => to_slv(opcode_type, 16#08#),
      3249 => to_slv(opcode_type, 16#07#),
      3250 => to_slv(opcode_type, 16#0F#),
      3251 => to_slv(opcode_type, 16#11#),
      3252 => to_slv(opcode_type, 16#08#),
      3253 => to_slv(opcode_type, 16#10#),
      3254 => to_slv(opcode_type, 16#59#),
      3255 => to_slv(opcode_type, 16#07#),
      3256 => to_slv(opcode_type, 16#08#),
      3257 => to_slv(opcode_type, 16#0E#),
      3258 => to_slv(opcode_type, 16#0B#),
      3259 => to_slv(opcode_type, 16#07#),
      3260 => to_slv(opcode_type, 16#0C#),
      3261 => to_slv(opcode_type, 16#0D#),
      3262 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#08#),
      3265 => to_slv(opcode_type, 16#07#),
      3266 => to_slv(opcode_type, 16#09#),
      3267 => to_slv(opcode_type, 16#02#),
      3268 => to_slv(opcode_type, 16#E2#),
      3269 => to_slv(opcode_type, 16#09#),
      3270 => to_slv(opcode_type, 16#0B#),
      3271 => to_slv(opcode_type, 16#0C#),
      3272 => to_slv(opcode_type, 16#06#),
      3273 => to_slv(opcode_type, 16#07#),
      3274 => to_slv(opcode_type, 16#10#),
      3275 => to_slv(opcode_type, 16#0C#),
      3276 => to_slv(opcode_type, 16#06#),
      3277 => to_slv(opcode_type, 16#0A#),
      3278 => to_slv(opcode_type, 16#0A#),
      3279 => to_slv(opcode_type, 16#07#),
      3280 => to_slv(opcode_type, 16#07#),
      3281 => to_slv(opcode_type, 16#09#),
      3282 => to_slv(opcode_type, 16#0E#),
      3283 => to_slv(opcode_type, 16#10#),
      3284 => to_slv(opcode_type, 16#08#),
      3285 => to_slv(opcode_type, 16#0E#),
      3286 => to_slv(opcode_type, 16#0C#),
      3287 => to_slv(opcode_type, 16#08#),
      3288 => to_slv(opcode_type, 16#06#),
      3289 => to_slv(opcode_type, 16#88#),
      3290 => to_slv(opcode_type, 16#A6#),
      3291 => to_slv(opcode_type, 16#06#),
      3292 => to_slv(opcode_type, 16#10#),
      3293 => to_slv(opcode_type, 16#0E#),
      3294 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#06#),
      3297 => to_slv(opcode_type, 16#09#),
      3298 => to_slv(opcode_type, 16#09#),
      3299 => to_slv(opcode_type, 16#07#),
      3300 => to_slv(opcode_type, 16#0F#),
      3301 => to_slv(opcode_type, 16#0C#),
      3302 => to_slv(opcode_type, 16#05#),
      3303 => to_slv(opcode_type, 16#84#),
      3304 => to_slv(opcode_type, 16#06#),
      3305 => to_slv(opcode_type, 16#09#),
      3306 => to_slv(opcode_type, 16#0B#),
      3307 => to_slv(opcode_type, 16#0D#),
      3308 => to_slv(opcode_type, 16#06#),
      3309 => to_slv(opcode_type, 16#10#),
      3310 => to_slv(opcode_type, 16#0C#),
      3311 => to_slv(opcode_type, 16#06#),
      3312 => to_slv(opcode_type, 16#09#),
      3313 => to_slv(opcode_type, 16#07#),
      3314 => to_slv(opcode_type, 16#B6#),
      3315 => to_slv(opcode_type, 16#11#),
      3316 => to_slv(opcode_type, 16#07#),
      3317 => to_slv(opcode_type, 16#11#),
      3318 => to_slv(opcode_type, 16#0F#),
      3319 => to_slv(opcode_type, 16#06#),
      3320 => to_slv(opcode_type, 16#06#),
      3321 => to_slv(opcode_type, 16#EB#),
      3322 => to_slv(opcode_type, 16#10#),
      3323 => to_slv(opcode_type, 16#06#),
      3324 => to_slv(opcode_type, 16#0F#),
      3325 => to_slv(opcode_type, 16#10#),
      3326 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#06#),
      3329 => to_slv(opcode_type, 16#07#),
      3330 => to_slv(opcode_type, 16#08#),
      3331 => to_slv(opcode_type, 16#02#),
      3332 => to_slv(opcode_type, 16#0B#),
      3333 => to_slv(opcode_type, 16#09#),
      3334 => to_slv(opcode_type, 16#0A#),
      3335 => to_slv(opcode_type, 16#0A#),
      3336 => to_slv(opcode_type, 16#08#),
      3337 => to_slv(opcode_type, 16#06#),
      3338 => to_slv(opcode_type, 16#0C#),
      3339 => to_slv(opcode_type, 16#7B#),
      3340 => to_slv(opcode_type, 16#07#),
      3341 => to_slv(opcode_type, 16#0C#),
      3342 => to_slv(opcode_type, 16#0F#),
      3343 => to_slv(opcode_type, 16#07#),
      3344 => to_slv(opcode_type, 16#06#),
      3345 => to_slv(opcode_type, 16#07#),
      3346 => to_slv(opcode_type, 16#0B#),
      3347 => to_slv(opcode_type, 16#0C#),
      3348 => to_slv(opcode_type, 16#08#),
      3349 => to_slv(opcode_type, 16#73#),
      3350 => to_slv(opcode_type, 16#0C#),
      3351 => to_slv(opcode_type, 16#07#),
      3352 => to_slv(opcode_type, 16#09#),
      3353 => to_slv(opcode_type, 16#0C#),
      3354 => to_slv(opcode_type, 16#0A#),
      3355 => to_slv(opcode_type, 16#07#),
      3356 => to_slv(opcode_type, 16#0E#),
      3357 => to_slv(opcode_type, 16#0B#),
      3358 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#08#),
      3361 => to_slv(opcode_type, 16#06#),
      3362 => to_slv(opcode_type, 16#06#),
      3363 => to_slv(opcode_type, 16#04#),
      3364 => to_slv(opcode_type, 16#0E#),
      3365 => to_slv(opcode_type, 16#07#),
      3366 => to_slv(opcode_type, 16#0F#),
      3367 => to_slv(opcode_type, 16#0C#),
      3368 => to_slv(opcode_type, 16#08#),
      3369 => to_slv(opcode_type, 16#08#),
      3370 => to_slv(opcode_type, 16#10#),
      3371 => to_slv(opcode_type, 16#0D#),
      3372 => to_slv(opcode_type, 16#06#),
      3373 => to_slv(opcode_type, 16#25#),
      3374 => to_slv(opcode_type, 16#10#),
      3375 => to_slv(opcode_type, 16#09#),
      3376 => to_slv(opcode_type, 16#09#),
      3377 => to_slv(opcode_type, 16#09#),
      3378 => to_slv(opcode_type, 16#0E#),
      3379 => to_slv(opcode_type, 16#10#),
      3380 => to_slv(opcode_type, 16#07#),
      3381 => to_slv(opcode_type, 16#0A#),
      3382 => to_slv(opcode_type, 16#0D#),
      3383 => to_slv(opcode_type, 16#08#),
      3384 => to_slv(opcode_type, 16#06#),
      3385 => to_slv(opcode_type, 16#11#),
      3386 => to_slv(opcode_type, 16#0A#),
      3387 => to_slv(opcode_type, 16#06#),
      3388 => to_slv(opcode_type, 16#0E#),
      3389 => to_slv(opcode_type, 16#0A#),
      3390 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#06#),
      3393 => to_slv(opcode_type, 16#07#),
      3394 => to_slv(opcode_type, 16#09#),
      3395 => to_slv(opcode_type, 16#04#),
      3396 => to_slv(opcode_type, 16#0B#),
      3397 => to_slv(opcode_type, 16#08#),
      3398 => to_slv(opcode_type, 16#0C#),
      3399 => to_slv(opcode_type, 16#30#),
      3400 => to_slv(opcode_type, 16#08#),
      3401 => to_slv(opcode_type, 16#09#),
      3402 => to_slv(opcode_type, 16#0F#),
      3403 => to_slv(opcode_type, 16#0A#),
      3404 => to_slv(opcode_type, 16#06#),
      3405 => to_slv(opcode_type, 16#0A#),
      3406 => to_slv(opcode_type, 16#0C#),
      3407 => to_slv(opcode_type, 16#06#),
      3408 => to_slv(opcode_type, 16#07#),
      3409 => to_slv(opcode_type, 16#09#),
      3410 => to_slv(opcode_type, 16#0B#),
      3411 => to_slv(opcode_type, 16#0F#),
      3412 => to_slv(opcode_type, 16#07#),
      3413 => to_slv(opcode_type, 16#89#),
      3414 => to_slv(opcode_type, 16#0E#),
      3415 => to_slv(opcode_type, 16#08#),
      3416 => to_slv(opcode_type, 16#07#),
      3417 => to_slv(opcode_type, 16#10#),
      3418 => to_slv(opcode_type, 16#11#),
      3419 => to_slv(opcode_type, 16#06#),
      3420 => to_slv(opcode_type, 16#0C#),
      3421 => to_slv(opcode_type, 16#10#),
      3422 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#08#),
      3425 => to_slv(opcode_type, 16#06#),
      3426 => to_slv(opcode_type, 16#06#),
      3427 => to_slv(opcode_type, 16#05#),
      3428 => to_slv(opcode_type, 16#0F#),
      3429 => to_slv(opcode_type, 16#09#),
      3430 => to_slv(opcode_type, 16#0B#),
      3431 => to_slv(opcode_type, 16#0E#),
      3432 => to_slv(opcode_type, 16#09#),
      3433 => to_slv(opcode_type, 16#06#),
      3434 => to_slv(opcode_type, 16#0E#),
      3435 => to_slv(opcode_type, 16#0C#),
      3436 => to_slv(opcode_type, 16#07#),
      3437 => to_slv(opcode_type, 16#11#),
      3438 => to_slv(opcode_type, 16#0E#),
      3439 => to_slv(opcode_type, 16#07#),
      3440 => to_slv(opcode_type, 16#07#),
      3441 => to_slv(opcode_type, 16#07#),
      3442 => to_slv(opcode_type, 16#0C#),
      3443 => to_slv(opcode_type, 16#0C#),
      3444 => to_slv(opcode_type, 16#09#),
      3445 => to_slv(opcode_type, 16#10#),
      3446 => to_slv(opcode_type, 16#0D#),
      3447 => to_slv(opcode_type, 16#08#),
      3448 => to_slv(opcode_type, 16#09#),
      3449 => to_slv(opcode_type, 16#0E#),
      3450 => to_slv(opcode_type, 16#0C#),
      3451 => to_slv(opcode_type, 16#07#),
      3452 => to_slv(opcode_type, 16#0F#),
      3453 => to_slv(opcode_type, 16#0A#),
      3454 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#07#),
      3457 => to_slv(opcode_type, 16#08#),
      3458 => to_slv(opcode_type, 16#08#),
      3459 => to_slv(opcode_type, 16#01#),
      3460 => to_slv(opcode_type, 16#11#),
      3461 => to_slv(opcode_type, 16#09#),
      3462 => to_slv(opcode_type, 16#0E#),
      3463 => to_slv(opcode_type, 16#0E#),
      3464 => to_slv(opcode_type, 16#06#),
      3465 => to_slv(opcode_type, 16#07#),
      3466 => to_slv(opcode_type, 16#0B#),
      3467 => to_slv(opcode_type, 16#70#),
      3468 => to_slv(opcode_type, 16#06#),
      3469 => to_slv(opcode_type, 16#0E#),
      3470 => to_slv(opcode_type, 16#0A#),
      3471 => to_slv(opcode_type, 16#09#),
      3472 => to_slv(opcode_type, 16#08#),
      3473 => to_slv(opcode_type, 16#09#),
      3474 => to_slv(opcode_type, 16#0E#),
      3475 => to_slv(opcode_type, 16#0F#),
      3476 => to_slv(opcode_type, 16#08#),
      3477 => to_slv(opcode_type, 16#0F#),
      3478 => to_slv(opcode_type, 16#0D#),
      3479 => to_slv(opcode_type, 16#07#),
      3480 => to_slv(opcode_type, 16#06#),
      3481 => to_slv(opcode_type, 16#0F#),
      3482 => to_slv(opcode_type, 16#11#),
      3483 => to_slv(opcode_type, 16#06#),
      3484 => to_slv(opcode_type, 16#0B#),
      3485 => to_slv(opcode_type, 16#0E#),
      3486 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#08#),
      3489 => to_slv(opcode_type, 16#06#),
      3490 => to_slv(opcode_type, 16#09#),
      3491 => to_slv(opcode_type, 16#06#),
      3492 => to_slv(opcode_type, 16#19#),
      3493 => to_slv(opcode_type, 16#9D#),
      3494 => to_slv(opcode_type, 16#09#),
      3495 => to_slv(opcode_type, 16#0B#),
      3496 => to_slv(opcode_type, 16#0B#),
      3497 => to_slv(opcode_type, 16#09#),
      3498 => to_slv(opcode_type, 16#04#),
      3499 => to_slv(opcode_type, 16#0F#),
      3500 => to_slv(opcode_type, 16#09#),
      3501 => to_slv(opcode_type, 16#97#),
      3502 => to_slv(opcode_type, 16#0C#),
      3503 => to_slv(opcode_type, 16#08#),
      3504 => to_slv(opcode_type, 16#09#),
      3505 => to_slv(opcode_type, 16#08#),
      3506 => to_slv(opcode_type, 16#10#),
      3507 => to_slv(opcode_type, 16#0C#),
      3508 => to_slv(opcode_type, 16#06#),
      3509 => to_slv(opcode_type, 16#10#),
      3510 => to_slv(opcode_type, 16#11#),
      3511 => to_slv(opcode_type, 16#06#),
      3512 => to_slv(opcode_type, 16#06#),
      3513 => to_slv(opcode_type, 16#0C#),
      3514 => to_slv(opcode_type, 16#0B#),
      3515 => to_slv(opcode_type, 16#08#),
      3516 => to_slv(opcode_type, 16#0B#),
      3517 => to_slv(opcode_type, 16#0B#),
      3518 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#06#),
      3521 => to_slv(opcode_type, 16#07#),
      3522 => to_slv(opcode_type, 16#09#),
      3523 => to_slv(opcode_type, 16#05#),
      3524 => to_slv(opcode_type, 16#0D#),
      3525 => to_slv(opcode_type, 16#08#),
      3526 => to_slv(opcode_type, 16#0D#),
      3527 => to_slv(opcode_type, 16#0F#),
      3528 => to_slv(opcode_type, 16#06#),
      3529 => to_slv(opcode_type, 16#09#),
      3530 => to_slv(opcode_type, 16#0B#),
      3531 => to_slv(opcode_type, 16#10#),
      3532 => to_slv(opcode_type, 16#09#),
      3533 => to_slv(opcode_type, 16#10#),
      3534 => to_slv(opcode_type, 16#11#),
      3535 => to_slv(opcode_type, 16#08#),
      3536 => to_slv(opcode_type, 16#08#),
      3537 => to_slv(opcode_type, 16#06#),
      3538 => to_slv(opcode_type, 16#0A#),
      3539 => to_slv(opcode_type, 16#11#),
      3540 => to_slv(opcode_type, 16#07#),
      3541 => to_slv(opcode_type, 16#0D#),
      3542 => to_slv(opcode_type, 16#0D#),
      3543 => to_slv(opcode_type, 16#08#),
      3544 => to_slv(opcode_type, 16#09#),
      3545 => to_slv(opcode_type, 16#11#),
      3546 => to_slv(opcode_type, 16#A3#),
      3547 => to_slv(opcode_type, 16#09#),
      3548 => to_slv(opcode_type, 16#0D#),
      3549 => to_slv(opcode_type, 16#0C#),
      3550 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#06#),
      3553 => to_slv(opcode_type, 16#09#),
      3554 => to_slv(opcode_type, 16#07#),
      3555 => to_slv(opcode_type, 16#09#),
      3556 => to_slv(opcode_type, 16#11#),
      3557 => to_slv(opcode_type, 16#0A#),
      3558 => to_slv(opcode_type, 16#06#),
      3559 => to_slv(opcode_type, 16#0D#),
      3560 => to_slv(opcode_type, 16#10#),
      3561 => to_slv(opcode_type, 16#08#),
      3562 => to_slv(opcode_type, 16#07#),
      3563 => to_slv(opcode_type, 16#0D#),
      3564 => to_slv(opcode_type, 16#0A#),
      3565 => to_slv(opcode_type, 16#02#),
      3566 => to_slv(opcode_type, 16#0E#),
      3567 => to_slv(opcode_type, 16#06#),
      3568 => to_slv(opcode_type, 16#09#),
      3569 => to_slv(opcode_type, 16#09#),
      3570 => to_slv(opcode_type, 16#B6#),
      3571 => to_slv(opcode_type, 16#0A#),
      3572 => to_slv(opcode_type, 16#08#),
      3573 => to_slv(opcode_type, 16#43#),
      3574 => to_slv(opcode_type, 16#0F#),
      3575 => to_slv(opcode_type, 16#09#),
      3576 => to_slv(opcode_type, 16#08#),
      3577 => to_slv(opcode_type, 16#10#),
      3578 => to_slv(opcode_type, 16#0B#),
      3579 => to_slv(opcode_type, 16#08#),
      3580 => to_slv(opcode_type, 16#0C#),
      3581 => to_slv(opcode_type, 16#0B#),
      3582 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#06#),
      3585 => to_slv(opcode_type, 16#06#),
      3586 => to_slv(opcode_type, 16#08#),
      3587 => to_slv(opcode_type, 16#07#),
      3588 => to_slv(opcode_type, 16#0D#),
      3589 => to_slv(opcode_type, 16#11#),
      3590 => to_slv(opcode_type, 16#06#),
      3591 => to_slv(opcode_type, 16#10#),
      3592 => to_slv(opcode_type, 16#10#),
      3593 => to_slv(opcode_type, 16#08#),
      3594 => to_slv(opcode_type, 16#01#),
      3595 => to_slv(opcode_type, 16#0A#),
      3596 => to_slv(opcode_type, 16#06#),
      3597 => to_slv(opcode_type, 16#10#),
      3598 => to_slv(opcode_type, 16#11#),
      3599 => to_slv(opcode_type, 16#06#),
      3600 => to_slv(opcode_type, 16#09#),
      3601 => to_slv(opcode_type, 16#06#),
      3602 => to_slv(opcode_type, 16#0A#),
      3603 => to_slv(opcode_type, 16#0C#),
      3604 => to_slv(opcode_type, 16#08#),
      3605 => to_slv(opcode_type, 16#0A#),
      3606 => to_slv(opcode_type, 16#0F#),
      3607 => to_slv(opcode_type, 16#08#),
      3608 => to_slv(opcode_type, 16#06#),
      3609 => to_slv(opcode_type, 16#85#),
      3610 => to_slv(opcode_type, 16#0A#),
      3611 => to_slv(opcode_type, 16#09#),
      3612 => to_slv(opcode_type, 16#10#),
      3613 => to_slv(opcode_type, 16#0C#),
      3614 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#09#),
      3617 => to_slv(opcode_type, 16#08#),
      3618 => to_slv(opcode_type, 16#09#),
      3619 => to_slv(opcode_type, 16#05#),
      3620 => to_slv(opcode_type, 16#10#),
      3621 => to_slv(opcode_type, 16#06#),
      3622 => to_slv(opcode_type, 16#D2#),
      3623 => to_slv(opcode_type, 16#0A#),
      3624 => to_slv(opcode_type, 16#07#),
      3625 => to_slv(opcode_type, 16#06#),
      3626 => to_slv(opcode_type, 16#11#),
      3627 => to_slv(opcode_type, 16#0A#),
      3628 => to_slv(opcode_type, 16#06#),
      3629 => to_slv(opcode_type, 16#0F#),
      3630 => to_slv(opcode_type, 16#11#),
      3631 => to_slv(opcode_type, 16#07#),
      3632 => to_slv(opcode_type, 16#07#),
      3633 => to_slv(opcode_type, 16#09#),
      3634 => to_slv(opcode_type, 16#0F#),
      3635 => to_slv(opcode_type, 16#0A#),
      3636 => to_slv(opcode_type, 16#06#),
      3637 => to_slv(opcode_type, 16#0B#),
      3638 => to_slv(opcode_type, 16#0F#),
      3639 => to_slv(opcode_type, 16#07#),
      3640 => to_slv(opcode_type, 16#07#),
      3641 => to_slv(opcode_type, 16#11#),
      3642 => to_slv(opcode_type, 16#0C#),
      3643 => to_slv(opcode_type, 16#09#),
      3644 => to_slv(opcode_type, 16#0B#),
      3645 => to_slv(opcode_type, 16#0A#),
      3646 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#06#),
      3649 => to_slv(opcode_type, 16#08#),
      3650 => to_slv(opcode_type, 16#06#),
      3651 => to_slv(opcode_type, 16#07#),
      3652 => to_slv(opcode_type, 16#0C#),
      3653 => to_slv(opcode_type, 16#0B#),
      3654 => to_slv(opcode_type, 16#06#),
      3655 => to_slv(opcode_type, 16#0C#),
      3656 => to_slv(opcode_type, 16#0C#),
      3657 => to_slv(opcode_type, 16#06#),
      3658 => to_slv(opcode_type, 16#06#),
      3659 => to_slv(opcode_type, 16#0B#),
      3660 => to_slv(opcode_type, 16#0D#),
      3661 => to_slv(opcode_type, 16#07#),
      3662 => to_slv(opcode_type, 16#0A#),
      3663 => to_slv(opcode_type, 16#0D#),
      3664 => to_slv(opcode_type, 16#08#),
      3665 => to_slv(opcode_type, 16#07#),
      3666 => to_slv(opcode_type, 16#06#),
      3667 => to_slv(opcode_type, 16#0D#),
      3668 => to_slv(opcode_type, 16#0B#),
      3669 => to_slv(opcode_type, 16#09#),
      3670 => to_slv(opcode_type, 16#0A#),
      3671 => to_slv(opcode_type, 16#F5#),
      3672 => to_slv(opcode_type, 16#06#),
      3673 => to_slv(opcode_type, 16#08#),
      3674 => to_slv(opcode_type, 16#EC#),
      3675 => to_slv(opcode_type, 16#10#),
      3676 => to_slv(opcode_type, 16#02#),
      3677 => to_slv(opcode_type, 16#0A#),
      3678 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#09#),
      3681 => to_slv(opcode_type, 16#07#),
      3682 => to_slv(opcode_type, 16#08#),
      3683 => to_slv(opcode_type, 16#05#),
      3684 => to_slv(opcode_type, 16#10#),
      3685 => to_slv(opcode_type, 16#09#),
      3686 => to_slv(opcode_type, 16#10#),
      3687 => to_slv(opcode_type, 16#34#),
      3688 => to_slv(opcode_type, 16#08#),
      3689 => to_slv(opcode_type, 16#09#),
      3690 => to_slv(opcode_type, 16#0E#),
      3691 => to_slv(opcode_type, 16#0D#),
      3692 => to_slv(opcode_type, 16#06#),
      3693 => to_slv(opcode_type, 16#0D#),
      3694 => to_slv(opcode_type, 16#0B#),
      3695 => to_slv(opcode_type, 16#07#),
      3696 => to_slv(opcode_type, 16#09#),
      3697 => to_slv(opcode_type, 16#07#),
      3698 => to_slv(opcode_type, 16#44#),
      3699 => to_slv(opcode_type, 16#11#),
      3700 => to_slv(opcode_type, 16#08#),
      3701 => to_slv(opcode_type, 16#0E#),
      3702 => to_slv(opcode_type, 16#0C#),
      3703 => to_slv(opcode_type, 16#08#),
      3704 => to_slv(opcode_type, 16#06#),
      3705 => to_slv(opcode_type, 16#0D#),
      3706 => to_slv(opcode_type, 16#0D#),
      3707 => to_slv(opcode_type, 16#08#),
      3708 => to_slv(opcode_type, 16#0D#),
      3709 => to_slv(opcode_type, 16#10#),
      3710 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#06#),
      3713 => to_slv(opcode_type, 16#09#),
      3714 => to_slv(opcode_type, 16#09#),
      3715 => to_slv(opcode_type, 16#04#),
      3716 => to_slv(opcode_type, 16#11#),
      3717 => to_slv(opcode_type, 16#07#),
      3718 => to_slv(opcode_type, 16#0C#),
      3719 => to_slv(opcode_type, 16#0B#),
      3720 => to_slv(opcode_type, 16#08#),
      3721 => to_slv(opcode_type, 16#08#),
      3722 => to_slv(opcode_type, 16#0D#),
      3723 => to_slv(opcode_type, 16#A8#),
      3724 => to_slv(opcode_type, 16#09#),
      3725 => to_slv(opcode_type, 16#0C#),
      3726 => to_slv(opcode_type, 16#0D#),
      3727 => to_slv(opcode_type, 16#09#),
      3728 => to_slv(opcode_type, 16#08#),
      3729 => to_slv(opcode_type, 16#06#),
      3730 => to_slv(opcode_type, 16#0F#),
      3731 => to_slv(opcode_type, 16#74#),
      3732 => to_slv(opcode_type, 16#09#),
      3733 => to_slv(opcode_type, 16#0F#),
      3734 => to_slv(opcode_type, 16#0D#),
      3735 => to_slv(opcode_type, 16#09#),
      3736 => to_slv(opcode_type, 16#08#),
      3737 => to_slv(opcode_type, 16#0B#),
      3738 => to_slv(opcode_type, 16#0E#),
      3739 => to_slv(opcode_type, 16#07#),
      3740 => to_slv(opcode_type, 16#0F#),
      3741 => to_slv(opcode_type, 16#0A#),
      3742 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#06#),
      3745 => to_slv(opcode_type, 16#07#),
      3746 => to_slv(opcode_type, 16#07#),
      3747 => to_slv(opcode_type, 16#04#),
      3748 => to_slv(opcode_type, 16#10#),
      3749 => to_slv(opcode_type, 16#06#),
      3750 => to_slv(opcode_type, 16#0A#),
      3751 => to_slv(opcode_type, 16#10#),
      3752 => to_slv(opcode_type, 16#08#),
      3753 => to_slv(opcode_type, 16#06#),
      3754 => to_slv(opcode_type, 16#E3#),
      3755 => to_slv(opcode_type, 16#0C#),
      3756 => to_slv(opcode_type, 16#06#),
      3757 => to_slv(opcode_type, 16#0A#),
      3758 => to_slv(opcode_type, 16#0A#),
      3759 => to_slv(opcode_type, 16#06#),
      3760 => to_slv(opcode_type, 16#09#),
      3761 => to_slv(opcode_type, 16#08#),
      3762 => to_slv(opcode_type, 16#10#),
      3763 => to_slv(opcode_type, 16#0B#),
      3764 => to_slv(opcode_type, 16#09#),
      3765 => to_slv(opcode_type, 16#0C#),
      3766 => to_slv(opcode_type, 16#0A#),
      3767 => to_slv(opcode_type, 16#06#),
      3768 => to_slv(opcode_type, 16#08#),
      3769 => to_slv(opcode_type, 16#CB#),
      3770 => to_slv(opcode_type, 16#0D#),
      3771 => to_slv(opcode_type, 16#08#),
      3772 => to_slv(opcode_type, 16#10#),
      3773 => to_slv(opcode_type, 16#0C#),
      3774 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#09#),
      3777 => to_slv(opcode_type, 16#07#),
      3778 => to_slv(opcode_type, 16#08#),
      3779 => to_slv(opcode_type, 16#02#),
      3780 => to_slv(opcode_type, 16#0A#),
      3781 => to_slv(opcode_type, 16#07#),
      3782 => to_slv(opcode_type, 16#11#),
      3783 => to_slv(opcode_type, 16#0B#),
      3784 => to_slv(opcode_type, 16#07#),
      3785 => to_slv(opcode_type, 16#09#),
      3786 => to_slv(opcode_type, 16#0A#),
      3787 => to_slv(opcode_type, 16#0C#),
      3788 => to_slv(opcode_type, 16#06#),
      3789 => to_slv(opcode_type, 16#10#),
      3790 => to_slv(opcode_type, 16#0B#),
      3791 => to_slv(opcode_type, 16#08#),
      3792 => to_slv(opcode_type, 16#06#),
      3793 => to_slv(opcode_type, 16#09#),
      3794 => to_slv(opcode_type, 16#0D#),
      3795 => to_slv(opcode_type, 16#0E#),
      3796 => to_slv(opcode_type, 16#07#),
      3797 => to_slv(opcode_type, 16#0B#),
      3798 => to_slv(opcode_type, 16#0B#),
      3799 => to_slv(opcode_type, 16#08#),
      3800 => to_slv(opcode_type, 16#06#),
      3801 => to_slv(opcode_type, 16#0B#),
      3802 => to_slv(opcode_type, 16#0C#),
      3803 => to_slv(opcode_type, 16#09#),
      3804 => to_slv(opcode_type, 16#0B#),
      3805 => to_slv(opcode_type, 16#0F#),
      3806 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#07#),
      3809 => to_slv(opcode_type, 16#07#),
      3810 => to_slv(opcode_type, 16#06#),
      3811 => to_slv(opcode_type, 16#08#),
      3812 => to_slv(opcode_type, 16#0F#),
      3813 => to_slv(opcode_type, 16#10#),
      3814 => to_slv(opcode_type, 16#08#),
      3815 => to_slv(opcode_type, 16#0F#),
      3816 => to_slv(opcode_type, 16#0A#),
      3817 => to_slv(opcode_type, 16#07#),
      3818 => to_slv(opcode_type, 16#07#),
      3819 => to_slv(opcode_type, 16#1F#),
      3820 => to_slv(opcode_type, 16#11#),
      3821 => to_slv(opcode_type, 16#09#),
      3822 => to_slv(opcode_type, 16#F9#),
      3823 => to_slv(opcode_type, 16#10#),
      3824 => to_slv(opcode_type, 16#07#),
      3825 => to_slv(opcode_type, 16#07#),
      3826 => to_slv(opcode_type, 16#01#),
      3827 => to_slv(opcode_type, 16#0A#),
      3828 => to_slv(opcode_type, 16#08#),
      3829 => to_slv(opcode_type, 16#0E#),
      3830 => to_slv(opcode_type, 16#0C#),
      3831 => to_slv(opcode_type, 16#07#),
      3832 => to_slv(opcode_type, 16#06#),
      3833 => to_slv(opcode_type, 16#0D#),
      3834 => to_slv(opcode_type, 16#0E#),
      3835 => to_slv(opcode_type, 16#07#),
      3836 => to_slv(opcode_type, 16#0B#),
      3837 => to_slv(opcode_type, 16#10#),
      3838 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#07#),
      3841 => to_slv(opcode_type, 16#08#),
      3842 => to_slv(opcode_type, 16#08#),
      3843 => to_slv(opcode_type, 16#06#),
      3844 => to_slv(opcode_type, 16#0B#),
      3845 => to_slv(opcode_type, 16#0D#),
      3846 => to_slv(opcode_type, 16#01#),
      3847 => to_slv(opcode_type, 16#0B#),
      3848 => to_slv(opcode_type, 16#06#),
      3849 => to_slv(opcode_type, 16#07#),
      3850 => to_slv(opcode_type, 16#0E#),
      3851 => to_slv(opcode_type, 16#10#),
      3852 => to_slv(opcode_type, 16#08#),
      3853 => to_slv(opcode_type, 16#10#),
      3854 => to_slv(opcode_type, 16#0E#),
      3855 => to_slv(opcode_type, 16#06#),
      3856 => to_slv(opcode_type, 16#06#),
      3857 => to_slv(opcode_type, 16#08#),
      3858 => to_slv(opcode_type, 16#F5#),
      3859 => to_slv(opcode_type, 16#0B#),
      3860 => to_slv(opcode_type, 16#07#),
      3861 => to_slv(opcode_type, 16#0C#),
      3862 => to_slv(opcode_type, 16#0A#),
      3863 => to_slv(opcode_type, 16#07#),
      3864 => to_slv(opcode_type, 16#07#),
      3865 => to_slv(opcode_type, 16#A6#),
      3866 => to_slv(opcode_type, 16#0A#),
      3867 => to_slv(opcode_type, 16#08#),
      3868 => to_slv(opcode_type, 16#0E#),
      3869 => to_slv(opcode_type, 16#0D#),
      3870 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#08#),
      3873 => to_slv(opcode_type, 16#07#),
      3874 => to_slv(opcode_type, 16#08#),
      3875 => to_slv(opcode_type, 16#07#),
      3876 => to_slv(opcode_type, 16#0C#),
      3877 => to_slv(opcode_type, 16#0C#),
      3878 => to_slv(opcode_type, 16#07#),
      3879 => to_slv(opcode_type, 16#CB#),
      3880 => to_slv(opcode_type, 16#0D#),
      3881 => to_slv(opcode_type, 16#06#),
      3882 => to_slv(opcode_type, 16#07#),
      3883 => to_slv(opcode_type, 16#11#),
      3884 => to_slv(opcode_type, 16#11#),
      3885 => to_slv(opcode_type, 16#03#),
      3886 => to_slv(opcode_type, 16#0A#),
      3887 => to_slv(opcode_type, 16#09#),
      3888 => to_slv(opcode_type, 16#09#),
      3889 => to_slv(opcode_type, 16#07#),
      3890 => to_slv(opcode_type, 16#0C#),
      3891 => to_slv(opcode_type, 16#0C#),
      3892 => to_slv(opcode_type, 16#09#),
      3893 => to_slv(opcode_type, 16#0B#),
      3894 => to_slv(opcode_type, 16#0D#),
      3895 => to_slv(opcode_type, 16#07#),
      3896 => to_slv(opcode_type, 16#08#),
      3897 => to_slv(opcode_type, 16#0B#),
      3898 => to_slv(opcode_type, 16#0C#),
      3899 => to_slv(opcode_type, 16#09#),
      3900 => to_slv(opcode_type, 16#0F#),
      3901 => to_slv(opcode_type, 16#0D#),
      3902 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#09#),
      3905 => to_slv(opcode_type, 16#06#),
      3906 => to_slv(opcode_type, 16#08#),
      3907 => to_slv(opcode_type, 16#04#),
      3908 => to_slv(opcode_type, 16#0F#),
      3909 => to_slv(opcode_type, 16#08#),
      3910 => to_slv(opcode_type, 16#11#),
      3911 => to_slv(opcode_type, 16#10#),
      3912 => to_slv(opcode_type, 16#06#),
      3913 => to_slv(opcode_type, 16#09#),
      3914 => to_slv(opcode_type, 16#62#),
      3915 => to_slv(opcode_type, 16#0D#),
      3916 => to_slv(opcode_type, 16#09#),
      3917 => to_slv(opcode_type, 16#0A#),
      3918 => to_slv(opcode_type, 16#0A#),
      3919 => to_slv(opcode_type, 16#07#),
      3920 => to_slv(opcode_type, 16#08#),
      3921 => to_slv(opcode_type, 16#09#),
      3922 => to_slv(opcode_type, 16#0A#),
      3923 => to_slv(opcode_type, 16#0A#),
      3924 => to_slv(opcode_type, 16#07#),
      3925 => to_slv(opcode_type, 16#10#),
      3926 => to_slv(opcode_type, 16#31#),
      3927 => to_slv(opcode_type, 16#07#),
      3928 => to_slv(opcode_type, 16#07#),
      3929 => to_slv(opcode_type, 16#10#),
      3930 => to_slv(opcode_type, 16#0B#),
      3931 => to_slv(opcode_type, 16#07#),
      3932 => to_slv(opcode_type, 16#11#),
      3933 => to_slv(opcode_type, 16#0A#),
      3934 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#07#),
      3937 => to_slv(opcode_type, 16#06#),
      3938 => to_slv(opcode_type, 16#06#),
      3939 => to_slv(opcode_type, 16#03#),
      3940 => to_slv(opcode_type, 16#0C#),
      3941 => to_slv(opcode_type, 16#09#),
      3942 => to_slv(opcode_type, 16#0C#),
      3943 => to_slv(opcode_type, 16#0B#),
      3944 => to_slv(opcode_type, 16#06#),
      3945 => to_slv(opcode_type, 16#06#),
      3946 => to_slv(opcode_type, 16#0A#),
      3947 => to_slv(opcode_type, 16#0A#),
      3948 => to_slv(opcode_type, 16#06#),
      3949 => to_slv(opcode_type, 16#11#),
      3950 => to_slv(opcode_type, 16#0E#),
      3951 => to_slv(opcode_type, 16#07#),
      3952 => to_slv(opcode_type, 16#08#),
      3953 => to_slv(opcode_type, 16#09#),
      3954 => to_slv(opcode_type, 16#0C#),
      3955 => to_slv(opcode_type, 16#0C#),
      3956 => to_slv(opcode_type, 16#07#),
      3957 => to_slv(opcode_type, 16#0B#),
      3958 => to_slv(opcode_type, 16#11#),
      3959 => to_slv(opcode_type, 16#08#),
      3960 => to_slv(opcode_type, 16#09#),
      3961 => to_slv(opcode_type, 16#0A#),
      3962 => to_slv(opcode_type, 16#0B#),
      3963 => to_slv(opcode_type, 16#07#),
      3964 => to_slv(opcode_type, 16#0A#),
      3965 => to_slv(opcode_type, 16#10#),
      3966 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#07#),
      3969 => to_slv(opcode_type, 16#06#),
      3970 => to_slv(opcode_type, 16#06#),
      3971 => to_slv(opcode_type, 16#08#),
      3972 => to_slv(opcode_type, 16#10#),
      3973 => to_slv(opcode_type, 16#0C#),
      3974 => to_slv(opcode_type, 16#09#),
      3975 => to_slv(opcode_type, 16#0B#),
      3976 => to_slv(opcode_type, 16#0E#),
      3977 => to_slv(opcode_type, 16#08#),
      3978 => to_slv(opcode_type, 16#02#),
      3979 => to_slv(opcode_type, 16#0B#),
      3980 => to_slv(opcode_type, 16#06#),
      3981 => to_slv(opcode_type, 16#0F#),
      3982 => to_slv(opcode_type, 16#0F#),
      3983 => to_slv(opcode_type, 16#07#),
      3984 => to_slv(opcode_type, 16#07#),
      3985 => to_slv(opcode_type, 16#07#),
      3986 => to_slv(opcode_type, 16#11#),
      3987 => to_slv(opcode_type, 16#0A#),
      3988 => to_slv(opcode_type, 16#08#),
      3989 => to_slv(opcode_type, 16#11#),
      3990 => to_slv(opcode_type, 16#0E#),
      3991 => to_slv(opcode_type, 16#07#),
      3992 => to_slv(opcode_type, 16#09#),
      3993 => to_slv(opcode_type, 16#0A#),
      3994 => to_slv(opcode_type, 16#10#),
      3995 => to_slv(opcode_type, 16#09#),
      3996 => to_slv(opcode_type, 16#0B#),
      3997 => to_slv(opcode_type, 16#10#),
      3998 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#07#),
      4001 => to_slv(opcode_type, 16#09#),
      4002 => to_slv(opcode_type, 16#06#),
      4003 => to_slv(opcode_type, 16#09#),
      4004 => to_slv(opcode_type, 16#0F#),
      4005 => to_slv(opcode_type, 16#0F#),
      4006 => to_slv(opcode_type, 16#04#),
      4007 => to_slv(opcode_type, 16#0C#),
      4008 => to_slv(opcode_type, 16#07#),
      4009 => to_slv(opcode_type, 16#08#),
      4010 => to_slv(opcode_type, 16#0E#),
      4011 => to_slv(opcode_type, 16#7B#),
      4012 => to_slv(opcode_type, 16#08#),
      4013 => to_slv(opcode_type, 16#1C#),
      4014 => to_slv(opcode_type, 16#0C#),
      4015 => to_slv(opcode_type, 16#07#),
      4016 => to_slv(opcode_type, 16#06#),
      4017 => to_slv(opcode_type, 16#08#),
      4018 => to_slv(opcode_type, 16#11#),
      4019 => to_slv(opcode_type, 16#D3#),
      4020 => to_slv(opcode_type, 16#08#),
      4021 => to_slv(opcode_type, 16#0E#),
      4022 => to_slv(opcode_type, 16#0C#),
      4023 => to_slv(opcode_type, 16#07#),
      4024 => to_slv(opcode_type, 16#07#),
      4025 => to_slv(opcode_type, 16#11#),
      4026 => to_slv(opcode_type, 16#0A#),
      4027 => to_slv(opcode_type, 16#06#),
      4028 => to_slv(opcode_type, 16#0B#),
      4029 => to_slv(opcode_type, 16#0C#),
      4030 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#08#),
      4033 => to_slv(opcode_type, 16#09#),
      4034 => to_slv(opcode_type, 16#08#),
      4035 => to_slv(opcode_type, 16#06#),
      4036 => to_slv(opcode_type, 16#0A#),
      4037 => to_slv(opcode_type, 16#11#),
      4038 => to_slv(opcode_type, 16#05#),
      4039 => to_slv(opcode_type, 16#0E#),
      4040 => to_slv(opcode_type, 16#09#),
      4041 => to_slv(opcode_type, 16#09#),
      4042 => to_slv(opcode_type, 16#11#),
      4043 => to_slv(opcode_type, 16#0D#),
      4044 => to_slv(opcode_type, 16#06#),
      4045 => to_slv(opcode_type, 16#32#),
      4046 => to_slv(opcode_type, 16#10#),
      4047 => to_slv(opcode_type, 16#09#),
      4048 => to_slv(opcode_type, 16#09#),
      4049 => to_slv(opcode_type, 16#09#),
      4050 => to_slv(opcode_type, 16#0D#),
      4051 => to_slv(opcode_type, 16#0C#),
      4052 => to_slv(opcode_type, 16#07#),
      4053 => to_slv(opcode_type, 16#0B#),
      4054 => to_slv(opcode_type, 16#0D#),
      4055 => to_slv(opcode_type, 16#09#),
      4056 => to_slv(opcode_type, 16#06#),
      4057 => to_slv(opcode_type, 16#0E#),
      4058 => to_slv(opcode_type, 16#0A#),
      4059 => to_slv(opcode_type, 16#09#),
      4060 => to_slv(opcode_type, 16#0E#),
      4061 => to_slv(opcode_type, 16#0A#),
      4062 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#08#),
      4065 => to_slv(opcode_type, 16#09#),
      4066 => to_slv(opcode_type, 16#09#),
      4067 => to_slv(opcode_type, 16#08#),
      4068 => to_slv(opcode_type, 16#0C#),
      4069 => to_slv(opcode_type, 16#0B#),
      4070 => to_slv(opcode_type, 16#02#),
      4071 => to_slv(opcode_type, 16#11#),
      4072 => to_slv(opcode_type, 16#09#),
      4073 => to_slv(opcode_type, 16#08#),
      4074 => to_slv(opcode_type, 16#0C#),
      4075 => to_slv(opcode_type, 16#10#),
      4076 => to_slv(opcode_type, 16#06#),
      4077 => to_slv(opcode_type, 16#0F#),
      4078 => to_slv(opcode_type, 16#10#),
      4079 => to_slv(opcode_type, 16#08#),
      4080 => to_slv(opcode_type, 16#09#),
      4081 => to_slv(opcode_type, 16#06#),
      4082 => to_slv(opcode_type, 16#B5#),
      4083 => to_slv(opcode_type, 16#0D#),
      4084 => to_slv(opcode_type, 16#07#),
      4085 => to_slv(opcode_type, 16#10#),
      4086 => to_slv(opcode_type, 16#0B#),
      4087 => to_slv(opcode_type, 16#08#),
      4088 => to_slv(opcode_type, 16#09#),
      4089 => to_slv(opcode_type, 16#0B#),
      4090 => to_slv(opcode_type, 16#0C#),
      4091 => to_slv(opcode_type, 16#09#),
      4092 => to_slv(opcode_type, 16#0D#),
      4093 => to_slv(opcode_type, 16#0B#),
      4094 to 4095 => (others => '0')
  ),

    -- Bin `31`...
    30 => (
      -- Program 0...
      0 => to_slv(opcode_type, 16#06#),
      1 => to_slv(opcode_type, 16#07#),
      2 => to_slv(opcode_type, 16#06#),
      3 => to_slv(opcode_type, 16#08#),
      4 => to_slv(opcode_type, 16#0E#),
      5 => to_slv(opcode_type, 16#0F#),
      6 => to_slv(opcode_type, 16#07#),
      7 => to_slv(opcode_type, 16#0C#),
      8 => to_slv(opcode_type, 16#0C#),
      9 => to_slv(opcode_type, 16#09#),
      10 => to_slv(opcode_type, 16#08#),
      11 => to_slv(opcode_type, 16#0B#),
      12 => to_slv(opcode_type, 16#0F#),
      13 => to_slv(opcode_type, 16#07#),
      14 => to_slv(opcode_type, 16#11#),
      15 => to_slv(opcode_type, 16#44#),
      16 => to_slv(opcode_type, 16#06#),
      17 => to_slv(opcode_type, 16#08#),
      18 => to_slv(opcode_type, 16#09#),
      19 => to_slv(opcode_type, 16#0E#),
      20 => to_slv(opcode_type, 16#0D#),
      21 => to_slv(opcode_type, 16#08#),
      22 => to_slv(opcode_type, 16#0E#),
      23 => to_slv(opcode_type, 16#0B#),
      24 => to_slv(opcode_type, 16#09#),
      25 => to_slv(opcode_type, 16#06#),
      26 => to_slv(opcode_type, 16#10#),
      27 => to_slv(opcode_type, 16#0B#),
      28 => to_slv(opcode_type, 16#08#),
      29 => to_slv(opcode_type, 16#11#),
      30 => to_slv(opcode_type, 16#0C#),
      31 to 31 => (others => '0'),

      -- Program 1...
      32 => to_slv(opcode_type, 16#08#),
      33 => to_slv(opcode_type, 16#08#),
      34 => to_slv(opcode_type, 16#07#),
      35 => to_slv(opcode_type, 16#06#),
      36 => to_slv(opcode_type, 16#0B#),
      37 => to_slv(opcode_type, 16#0E#),
      38 => to_slv(opcode_type, 16#06#),
      39 => to_slv(opcode_type, 16#0C#),
      40 => to_slv(opcode_type, 16#0E#),
      41 => to_slv(opcode_type, 16#08#),
      42 => to_slv(opcode_type, 16#08#),
      43 => to_slv(opcode_type, 16#0D#),
      44 => to_slv(opcode_type, 16#0B#),
      45 => to_slv(opcode_type, 16#07#),
      46 => to_slv(opcode_type, 16#0A#),
      47 => to_slv(opcode_type, 16#0D#),
      48 => to_slv(opcode_type, 16#06#),
      49 => to_slv(opcode_type, 16#09#),
      50 => to_slv(opcode_type, 16#06#),
      51 => to_slv(opcode_type, 16#0D#),
      52 => to_slv(opcode_type, 16#0C#),
      53 => to_slv(opcode_type, 16#07#),
      54 => to_slv(opcode_type, 16#0E#),
      55 => to_slv(opcode_type, 16#12#),
      56 => to_slv(opcode_type, 16#07#),
      57 => to_slv(opcode_type, 16#08#),
      58 => to_slv(opcode_type, 16#0D#),
      59 => to_slv(opcode_type, 16#31#),
      60 => to_slv(opcode_type, 16#06#),
      61 => to_slv(opcode_type, 16#0F#),
      62 => to_slv(opcode_type, 16#10#),
      63 to 63 => (others => '0'),

      -- Program 2...
      64 => to_slv(opcode_type, 16#06#),
      65 => to_slv(opcode_type, 16#07#),
      66 => to_slv(opcode_type, 16#06#),
      67 => to_slv(opcode_type, 16#06#),
      68 => to_slv(opcode_type, 16#0E#),
      69 => to_slv(opcode_type, 16#0B#),
      70 => to_slv(opcode_type, 16#06#),
      71 => to_slv(opcode_type, 16#0D#),
      72 => to_slv(opcode_type, 16#0B#),
      73 => to_slv(opcode_type, 16#06#),
      74 => to_slv(opcode_type, 16#06#),
      75 => to_slv(opcode_type, 16#0F#),
      76 => to_slv(opcode_type, 16#0C#),
      77 => to_slv(opcode_type, 16#06#),
      78 => to_slv(opcode_type, 16#0E#),
      79 => to_slv(opcode_type, 16#0D#),
      80 => to_slv(opcode_type, 16#09#),
      81 => to_slv(opcode_type, 16#08#),
      82 => to_slv(opcode_type, 16#08#),
      83 => to_slv(opcode_type, 16#0C#),
      84 => to_slv(opcode_type, 16#0F#),
      85 => to_slv(opcode_type, 16#07#),
      86 => to_slv(opcode_type, 16#10#),
      87 => to_slv(opcode_type, 16#0B#),
      88 => to_slv(opcode_type, 16#08#),
      89 => to_slv(opcode_type, 16#07#),
      90 => to_slv(opcode_type, 16#0F#),
      91 => to_slv(opcode_type, 16#0E#),
      92 => to_slv(opcode_type, 16#09#),
      93 => to_slv(opcode_type, 16#0D#),
      94 => to_slv(opcode_type, 16#10#),
      95 to 95 => (others => '0'),

      -- Program 3...
      96 => to_slv(opcode_type, 16#06#),
      97 => to_slv(opcode_type, 16#08#),
      98 => to_slv(opcode_type, 16#07#),
      99 => to_slv(opcode_type, 16#06#),
      100 => to_slv(opcode_type, 16#0A#),
      101 => to_slv(opcode_type, 16#0E#),
      102 => to_slv(opcode_type, 16#06#),
      103 => to_slv(opcode_type, 16#0F#),
      104 => to_slv(opcode_type, 16#0F#),
      105 => to_slv(opcode_type, 16#09#),
      106 => to_slv(opcode_type, 16#07#),
      107 => to_slv(opcode_type, 16#42#),
      108 => to_slv(opcode_type, 16#10#),
      109 => to_slv(opcode_type, 16#09#),
      110 => to_slv(opcode_type, 16#0F#),
      111 => to_slv(opcode_type, 16#0E#),
      112 => to_slv(opcode_type, 16#06#),
      113 => to_slv(opcode_type, 16#09#),
      114 => to_slv(opcode_type, 16#06#),
      115 => to_slv(opcode_type, 16#0C#),
      116 => to_slv(opcode_type, 16#0A#),
      117 => to_slv(opcode_type, 16#07#),
      118 => to_slv(opcode_type, 16#10#),
      119 => to_slv(opcode_type, 16#0F#),
      120 => to_slv(opcode_type, 16#06#),
      121 => to_slv(opcode_type, 16#08#),
      122 => to_slv(opcode_type, 16#F9#),
      123 => to_slv(opcode_type, 16#0F#),
      124 => to_slv(opcode_type, 16#09#),
      125 => to_slv(opcode_type, 16#1C#),
      126 => to_slv(opcode_type, 16#0C#),
      127 to 127 => (others => '0'),

      -- Program 4...
      128 => to_slv(opcode_type, 16#09#),
      129 => to_slv(opcode_type, 16#07#),
      130 => to_slv(opcode_type, 16#07#),
      131 => to_slv(opcode_type, 16#07#),
      132 => to_slv(opcode_type, 16#3C#),
      133 => to_slv(opcode_type, 16#0E#),
      134 => to_slv(opcode_type, 16#07#),
      135 => to_slv(opcode_type, 16#11#),
      136 => to_slv(opcode_type, 16#0C#),
      137 => to_slv(opcode_type, 16#06#),
      138 => to_slv(opcode_type, 16#09#),
      139 => to_slv(opcode_type, 16#11#),
      140 => to_slv(opcode_type, 16#0D#),
      141 => to_slv(opcode_type, 16#09#),
      142 => to_slv(opcode_type, 16#0C#),
      143 => to_slv(opcode_type, 16#0B#),
      144 => to_slv(opcode_type, 16#06#),
      145 => to_slv(opcode_type, 16#06#),
      146 => to_slv(opcode_type, 16#09#),
      147 => to_slv(opcode_type, 16#0B#),
      148 => to_slv(opcode_type, 16#0A#),
      149 => to_slv(opcode_type, 16#07#),
      150 => to_slv(opcode_type, 16#11#),
      151 => to_slv(opcode_type, 16#0A#),
      152 => to_slv(opcode_type, 16#08#),
      153 => to_slv(opcode_type, 16#08#),
      154 => to_slv(opcode_type, 16#0D#),
      155 => to_slv(opcode_type, 16#0F#),
      156 => to_slv(opcode_type, 16#07#),
      157 => to_slv(opcode_type, 16#0D#),
      158 => to_slv(opcode_type, 16#0A#),
      159 to 159 => (others => '0'),

      -- Program 5...
      160 => to_slv(opcode_type, 16#06#),
      161 => to_slv(opcode_type, 16#07#),
      162 => to_slv(opcode_type, 16#08#),
      163 => to_slv(opcode_type, 16#09#),
      164 => to_slv(opcode_type, 16#0E#),
      165 => to_slv(opcode_type, 16#0B#),
      166 => to_slv(opcode_type, 16#08#),
      167 => to_slv(opcode_type, 16#CB#),
      168 => to_slv(opcode_type, 16#11#),
      169 => to_slv(opcode_type, 16#08#),
      170 => to_slv(opcode_type, 16#07#),
      171 => to_slv(opcode_type, 16#11#),
      172 => to_slv(opcode_type, 16#0A#),
      173 => to_slv(opcode_type, 16#06#),
      174 => to_slv(opcode_type, 16#0D#),
      175 => to_slv(opcode_type, 16#0E#),
      176 => to_slv(opcode_type, 16#07#),
      177 => to_slv(opcode_type, 16#07#),
      178 => to_slv(opcode_type, 16#08#),
      179 => to_slv(opcode_type, 16#0F#),
      180 => to_slv(opcode_type, 16#0C#),
      181 => to_slv(opcode_type, 16#08#),
      182 => to_slv(opcode_type, 16#0A#),
      183 => to_slv(opcode_type, 16#0D#),
      184 => to_slv(opcode_type, 16#06#),
      185 => to_slv(opcode_type, 16#08#),
      186 => to_slv(opcode_type, 16#B3#),
      187 => to_slv(opcode_type, 16#10#),
      188 => to_slv(opcode_type, 16#07#),
      189 => to_slv(opcode_type, 16#0D#),
      190 => to_slv(opcode_type, 16#0A#),
      191 to 191 => (others => '0'),

      -- Program 6...
      192 => to_slv(opcode_type, 16#08#),
      193 => to_slv(opcode_type, 16#09#),
      194 => to_slv(opcode_type, 16#06#),
      195 => to_slv(opcode_type, 16#07#),
      196 => to_slv(opcode_type, 16#11#),
      197 => to_slv(opcode_type, 16#11#),
      198 => to_slv(opcode_type, 16#06#),
      199 => to_slv(opcode_type, 16#11#),
      200 => to_slv(opcode_type, 16#BF#),
      201 => to_slv(opcode_type, 16#06#),
      202 => to_slv(opcode_type, 16#08#),
      203 => to_slv(opcode_type, 16#0C#),
      204 => to_slv(opcode_type, 16#0F#),
      205 => to_slv(opcode_type, 16#09#),
      206 => to_slv(opcode_type, 16#8E#),
      207 => to_slv(opcode_type, 16#0A#),
      208 => to_slv(opcode_type, 16#06#),
      209 => to_slv(opcode_type, 16#06#),
      210 => to_slv(opcode_type, 16#06#),
      211 => to_slv(opcode_type, 16#0C#),
      212 => to_slv(opcode_type, 16#0A#),
      213 => to_slv(opcode_type, 16#06#),
      214 => to_slv(opcode_type, 16#0F#),
      215 => to_slv(opcode_type, 16#0C#),
      216 => to_slv(opcode_type, 16#06#),
      217 => to_slv(opcode_type, 16#09#),
      218 => to_slv(opcode_type, 16#0B#),
      219 => to_slv(opcode_type, 16#0D#),
      220 => to_slv(opcode_type, 16#09#),
      221 => to_slv(opcode_type, 16#0F#),
      222 => to_slv(opcode_type, 16#0F#),
      223 to 223 => (others => '0'),

      -- Program 7...
      224 => to_slv(opcode_type, 16#07#),
      225 => to_slv(opcode_type, 16#08#),
      226 => to_slv(opcode_type, 16#06#),
      227 => to_slv(opcode_type, 16#07#),
      228 => to_slv(opcode_type, 16#0A#),
      229 => to_slv(opcode_type, 16#D4#),
      230 => to_slv(opcode_type, 16#06#),
      231 => to_slv(opcode_type, 16#0C#),
      232 => to_slv(opcode_type, 16#0F#),
      233 => to_slv(opcode_type, 16#06#),
      234 => to_slv(opcode_type, 16#07#),
      235 => to_slv(opcode_type, 16#80#),
      236 => to_slv(opcode_type, 16#0C#),
      237 => to_slv(opcode_type, 16#06#),
      238 => to_slv(opcode_type, 16#7D#),
      239 => to_slv(opcode_type, 16#0C#),
      240 => to_slv(opcode_type, 16#06#),
      241 => to_slv(opcode_type, 16#07#),
      242 => to_slv(opcode_type, 16#09#),
      243 => to_slv(opcode_type, 16#0E#),
      244 => to_slv(opcode_type, 16#0C#),
      245 => to_slv(opcode_type, 16#08#),
      246 => to_slv(opcode_type, 16#0D#),
      247 => to_slv(opcode_type, 16#0E#),
      248 => to_slv(opcode_type, 16#07#),
      249 => to_slv(opcode_type, 16#06#),
      250 => to_slv(opcode_type, 16#0D#),
      251 => to_slv(opcode_type, 16#0E#),
      252 => to_slv(opcode_type, 16#09#),
      253 => to_slv(opcode_type, 16#0E#),
      254 => to_slv(opcode_type, 16#0F#),
      255 to 255 => (others => '0'),

      -- Program 8...
      256 => to_slv(opcode_type, 16#09#),
      257 => to_slv(opcode_type, 16#06#),
      258 => to_slv(opcode_type, 16#06#),
      259 => to_slv(opcode_type, 16#07#),
      260 => to_slv(opcode_type, 16#0B#),
      261 => to_slv(opcode_type, 16#10#),
      262 => to_slv(opcode_type, 16#06#),
      263 => to_slv(opcode_type, 16#0C#),
      264 => to_slv(opcode_type, 16#0B#),
      265 => to_slv(opcode_type, 16#09#),
      266 => to_slv(opcode_type, 16#09#),
      267 => to_slv(opcode_type, 16#10#),
      268 => to_slv(opcode_type, 16#0A#),
      269 => to_slv(opcode_type, 16#09#),
      270 => to_slv(opcode_type, 16#0D#),
      271 => to_slv(opcode_type, 16#0C#),
      272 => to_slv(opcode_type, 16#07#),
      273 => to_slv(opcode_type, 16#08#),
      274 => to_slv(opcode_type, 16#09#),
      275 => to_slv(opcode_type, 16#0F#),
      276 => to_slv(opcode_type, 16#0F#),
      277 => to_slv(opcode_type, 16#09#),
      278 => to_slv(opcode_type, 16#0C#),
      279 => to_slv(opcode_type, 16#0B#),
      280 => to_slv(opcode_type, 16#09#),
      281 => to_slv(opcode_type, 16#06#),
      282 => to_slv(opcode_type, 16#2F#),
      283 => to_slv(opcode_type, 16#11#),
      284 => to_slv(opcode_type, 16#08#),
      285 => to_slv(opcode_type, 16#0A#),
      286 => to_slv(opcode_type, 16#10#),
      287 to 287 => (others => '0'),

      -- Program 9...
      288 => to_slv(opcode_type, 16#07#),
      289 => to_slv(opcode_type, 16#06#),
      290 => to_slv(opcode_type, 16#07#),
      291 => to_slv(opcode_type, 16#08#),
      292 => to_slv(opcode_type, 16#0E#),
      293 => to_slv(opcode_type, 16#0E#),
      294 => to_slv(opcode_type, 16#09#),
      295 => to_slv(opcode_type, 16#0A#),
      296 => to_slv(opcode_type, 16#0B#),
      297 => to_slv(opcode_type, 16#08#),
      298 => to_slv(opcode_type, 16#09#),
      299 => to_slv(opcode_type, 16#0A#),
      300 => to_slv(opcode_type, 16#D5#),
      301 => to_slv(opcode_type, 16#08#),
      302 => to_slv(opcode_type, 16#0E#),
      303 => to_slv(opcode_type, 16#F1#),
      304 => to_slv(opcode_type, 16#08#),
      305 => to_slv(opcode_type, 16#07#),
      306 => to_slv(opcode_type, 16#06#),
      307 => to_slv(opcode_type, 16#0C#),
      308 => to_slv(opcode_type, 16#0D#),
      309 => to_slv(opcode_type, 16#08#),
      310 => to_slv(opcode_type, 16#0E#),
      311 => to_slv(opcode_type, 16#0F#),
      312 => to_slv(opcode_type, 16#09#),
      313 => to_slv(opcode_type, 16#07#),
      314 => to_slv(opcode_type, 16#0E#),
      315 => to_slv(opcode_type, 16#10#),
      316 => to_slv(opcode_type, 16#06#),
      317 => to_slv(opcode_type, 16#18#),
      318 => to_slv(opcode_type, 16#0A#),
      319 to 319 => (others => '0'),

      -- Program 10...
      320 => to_slv(opcode_type, 16#08#),
      321 => to_slv(opcode_type, 16#07#),
      322 => to_slv(opcode_type, 16#06#),
      323 => to_slv(opcode_type, 16#06#),
      324 => to_slv(opcode_type, 16#0F#),
      325 => to_slv(opcode_type, 16#11#),
      326 => to_slv(opcode_type, 16#08#),
      327 => to_slv(opcode_type, 16#18#),
      328 => to_slv(opcode_type, 16#0D#),
      329 => to_slv(opcode_type, 16#06#),
      330 => to_slv(opcode_type, 16#07#),
      331 => to_slv(opcode_type, 16#4C#),
      332 => to_slv(opcode_type, 16#0E#),
      333 => to_slv(opcode_type, 16#06#),
      334 => to_slv(opcode_type, 16#0A#),
      335 => to_slv(opcode_type, 16#0A#),
      336 => to_slv(opcode_type, 16#08#),
      337 => to_slv(opcode_type, 16#09#),
      338 => to_slv(opcode_type, 16#06#),
      339 => to_slv(opcode_type, 16#0B#),
      340 => to_slv(opcode_type, 16#0B#),
      341 => to_slv(opcode_type, 16#09#),
      342 => to_slv(opcode_type, 16#0A#),
      343 => to_slv(opcode_type, 16#0F#),
      344 => to_slv(opcode_type, 16#07#),
      345 => to_slv(opcode_type, 16#08#),
      346 => to_slv(opcode_type, 16#0A#),
      347 => to_slv(opcode_type, 16#0E#),
      348 => to_slv(opcode_type, 16#08#),
      349 => to_slv(opcode_type, 16#0A#),
      350 => to_slv(opcode_type, 16#10#),
      351 to 351 => (others => '0'),

      -- Program 11...
      352 => to_slv(opcode_type, 16#07#),
      353 => to_slv(opcode_type, 16#09#),
      354 => to_slv(opcode_type, 16#09#),
      355 => to_slv(opcode_type, 16#07#),
      356 => to_slv(opcode_type, 16#11#),
      357 => to_slv(opcode_type, 16#0A#),
      358 => to_slv(opcode_type, 16#09#),
      359 => to_slv(opcode_type, 16#0C#),
      360 => to_slv(opcode_type, 16#0B#),
      361 => to_slv(opcode_type, 16#06#),
      362 => to_slv(opcode_type, 16#07#),
      363 => to_slv(opcode_type, 16#0A#),
      364 => to_slv(opcode_type, 16#0B#),
      365 => to_slv(opcode_type, 16#08#),
      366 => to_slv(opcode_type, 16#10#),
      367 => to_slv(opcode_type, 16#21#),
      368 => to_slv(opcode_type, 16#07#),
      369 => to_slv(opcode_type, 16#08#),
      370 => to_slv(opcode_type, 16#09#),
      371 => to_slv(opcode_type, 16#0B#),
      372 => to_slv(opcode_type, 16#0D#),
      373 => to_slv(opcode_type, 16#07#),
      374 => to_slv(opcode_type, 16#11#),
      375 => to_slv(opcode_type, 16#0E#),
      376 => to_slv(opcode_type, 16#06#),
      377 => to_slv(opcode_type, 16#09#),
      378 => to_slv(opcode_type, 16#0A#),
      379 => to_slv(opcode_type, 16#0F#),
      380 => to_slv(opcode_type, 16#07#),
      381 => to_slv(opcode_type, 16#0F#),
      382 => to_slv(opcode_type, 16#0D#),
      383 to 383 => (others => '0'),

      -- Program 12...
      384 => to_slv(opcode_type, 16#09#),
      385 => to_slv(opcode_type, 16#06#),
      386 => to_slv(opcode_type, 16#07#),
      387 => to_slv(opcode_type, 16#08#),
      388 => to_slv(opcode_type, 16#0E#),
      389 => to_slv(opcode_type, 16#10#),
      390 => to_slv(opcode_type, 16#08#),
      391 => to_slv(opcode_type, 16#D7#),
      392 => to_slv(opcode_type, 16#F5#),
      393 => to_slv(opcode_type, 16#07#),
      394 => to_slv(opcode_type, 16#09#),
      395 => to_slv(opcode_type, 16#10#),
      396 => to_slv(opcode_type, 16#0A#),
      397 => to_slv(opcode_type, 16#06#),
      398 => to_slv(opcode_type, 16#0B#),
      399 => to_slv(opcode_type, 16#0D#),
      400 => to_slv(opcode_type, 16#07#),
      401 => to_slv(opcode_type, 16#09#),
      402 => to_slv(opcode_type, 16#07#),
      403 => to_slv(opcode_type, 16#11#),
      404 => to_slv(opcode_type, 16#10#),
      405 => to_slv(opcode_type, 16#07#),
      406 => to_slv(opcode_type, 16#0D#),
      407 => to_slv(opcode_type, 16#0E#),
      408 => to_slv(opcode_type, 16#08#),
      409 => to_slv(opcode_type, 16#09#),
      410 => to_slv(opcode_type, 16#11#),
      411 => to_slv(opcode_type, 16#0B#),
      412 => to_slv(opcode_type, 16#07#),
      413 => to_slv(opcode_type, 16#0D#),
      414 => to_slv(opcode_type, 16#0A#),
      415 to 415 => (others => '0'),

      -- Program 13...
      416 => to_slv(opcode_type, 16#06#),
      417 => to_slv(opcode_type, 16#08#),
      418 => to_slv(opcode_type, 16#07#),
      419 => to_slv(opcode_type, 16#09#),
      420 => to_slv(opcode_type, 16#0D#),
      421 => to_slv(opcode_type, 16#0B#),
      422 => to_slv(opcode_type, 16#09#),
      423 => to_slv(opcode_type, 16#11#),
      424 => to_slv(opcode_type, 16#11#),
      425 => to_slv(opcode_type, 16#07#),
      426 => to_slv(opcode_type, 16#06#),
      427 => to_slv(opcode_type, 16#0C#),
      428 => to_slv(opcode_type, 16#0C#),
      429 => to_slv(opcode_type, 16#07#),
      430 => to_slv(opcode_type, 16#0C#),
      431 => to_slv(opcode_type, 16#0F#),
      432 => to_slv(opcode_type, 16#06#),
      433 => to_slv(opcode_type, 16#08#),
      434 => to_slv(opcode_type, 16#06#),
      435 => to_slv(opcode_type, 16#11#),
      436 => to_slv(opcode_type, 16#25#),
      437 => to_slv(opcode_type, 16#09#),
      438 => to_slv(opcode_type, 16#0D#),
      439 => to_slv(opcode_type, 16#6D#),
      440 => to_slv(opcode_type, 16#08#),
      441 => to_slv(opcode_type, 16#07#),
      442 => to_slv(opcode_type, 16#10#),
      443 => to_slv(opcode_type, 16#F9#),
      444 => to_slv(opcode_type, 16#08#),
      445 => to_slv(opcode_type, 16#10#),
      446 => to_slv(opcode_type, 16#0A#),
      447 to 447 => (others => '0'),

      -- Program 14...
      448 => to_slv(opcode_type, 16#08#),
      449 => to_slv(opcode_type, 16#08#),
      450 => to_slv(opcode_type, 16#09#),
      451 => to_slv(opcode_type, 16#07#),
      452 => to_slv(opcode_type, 16#0B#),
      453 => to_slv(opcode_type, 16#0E#),
      454 => to_slv(opcode_type, 16#09#),
      455 => to_slv(opcode_type, 16#0B#),
      456 => to_slv(opcode_type, 16#0A#),
      457 => to_slv(opcode_type, 16#07#),
      458 => to_slv(opcode_type, 16#09#),
      459 => to_slv(opcode_type, 16#0F#),
      460 => to_slv(opcode_type, 16#0A#),
      461 => to_slv(opcode_type, 16#08#),
      462 => to_slv(opcode_type, 16#0E#),
      463 => to_slv(opcode_type, 16#0C#),
      464 => to_slv(opcode_type, 16#09#),
      465 => to_slv(opcode_type, 16#08#),
      466 => to_slv(opcode_type, 16#08#),
      467 => to_slv(opcode_type, 16#0B#),
      468 => to_slv(opcode_type, 16#0B#),
      469 => to_slv(opcode_type, 16#09#),
      470 => to_slv(opcode_type, 16#0A#),
      471 => to_slv(opcode_type, 16#0E#),
      472 => to_slv(opcode_type, 16#08#),
      473 => to_slv(opcode_type, 16#09#),
      474 => to_slv(opcode_type, 16#B4#),
      475 => to_slv(opcode_type, 16#11#),
      476 => to_slv(opcode_type, 16#06#),
      477 => to_slv(opcode_type, 16#0D#),
      478 => to_slv(opcode_type, 16#0C#),
      479 to 479 => (others => '0'),

      -- Program 15...
      480 => to_slv(opcode_type, 16#06#),
      481 => to_slv(opcode_type, 16#07#),
      482 => to_slv(opcode_type, 16#08#),
      483 => to_slv(opcode_type, 16#07#),
      484 => to_slv(opcode_type, 16#0C#),
      485 => to_slv(opcode_type, 16#D9#),
      486 => to_slv(opcode_type, 16#07#),
      487 => to_slv(opcode_type, 16#0A#),
      488 => to_slv(opcode_type, 16#0C#),
      489 => to_slv(opcode_type, 16#06#),
      490 => to_slv(opcode_type, 16#07#),
      491 => to_slv(opcode_type, 16#10#),
      492 => to_slv(opcode_type, 16#10#),
      493 => to_slv(opcode_type, 16#07#),
      494 => to_slv(opcode_type, 16#0B#),
      495 => to_slv(opcode_type, 16#0F#),
      496 => to_slv(opcode_type, 16#08#),
      497 => to_slv(opcode_type, 16#08#),
      498 => to_slv(opcode_type, 16#06#),
      499 => to_slv(opcode_type, 16#0D#),
      500 => to_slv(opcode_type, 16#0A#),
      501 => to_slv(opcode_type, 16#08#),
      502 => to_slv(opcode_type, 16#10#),
      503 => to_slv(opcode_type, 16#0D#),
      504 => to_slv(opcode_type, 16#09#),
      505 => to_slv(opcode_type, 16#07#),
      506 => to_slv(opcode_type, 16#0A#),
      507 => to_slv(opcode_type, 16#0D#),
      508 => to_slv(opcode_type, 16#08#),
      509 => to_slv(opcode_type, 16#0F#),
      510 => to_slv(opcode_type, 16#0C#),
      511 to 511 => (others => '0'),

      -- Program 16...
      512 => to_slv(opcode_type, 16#09#),
      513 => to_slv(opcode_type, 16#07#),
      514 => to_slv(opcode_type, 16#07#),
      515 => to_slv(opcode_type, 16#06#),
      516 => to_slv(opcode_type, 16#0C#),
      517 => to_slv(opcode_type, 16#0E#),
      518 => to_slv(opcode_type, 16#06#),
      519 => to_slv(opcode_type, 16#0C#),
      520 => to_slv(opcode_type, 16#10#),
      521 => to_slv(opcode_type, 16#06#),
      522 => to_slv(opcode_type, 16#08#),
      523 => to_slv(opcode_type, 16#0D#),
      524 => to_slv(opcode_type, 16#0D#),
      525 => to_slv(opcode_type, 16#06#),
      526 => to_slv(opcode_type, 16#0C#),
      527 => to_slv(opcode_type, 16#0F#),
      528 => to_slv(opcode_type, 16#07#),
      529 => to_slv(opcode_type, 16#09#),
      530 => to_slv(opcode_type, 16#06#),
      531 => to_slv(opcode_type, 16#0A#),
      532 => to_slv(opcode_type, 16#0C#),
      533 => to_slv(opcode_type, 16#08#),
      534 => to_slv(opcode_type, 16#0E#),
      535 => to_slv(opcode_type, 16#0B#),
      536 => to_slv(opcode_type, 16#07#),
      537 => to_slv(opcode_type, 16#06#),
      538 => to_slv(opcode_type, 16#94#),
      539 => to_slv(opcode_type, 16#0A#),
      540 => to_slv(opcode_type, 16#07#),
      541 => to_slv(opcode_type, 16#0B#),
      542 => to_slv(opcode_type, 16#2E#),
      543 to 543 => (others => '0'),

      -- Program 17...
      544 => to_slv(opcode_type, 16#09#),
      545 => to_slv(opcode_type, 16#06#),
      546 => to_slv(opcode_type, 16#08#),
      547 => to_slv(opcode_type, 16#07#),
      548 => to_slv(opcode_type, 16#0C#),
      549 => to_slv(opcode_type, 16#0E#),
      550 => to_slv(opcode_type, 16#09#),
      551 => to_slv(opcode_type, 16#9C#),
      552 => to_slv(opcode_type, 16#0F#),
      553 => to_slv(opcode_type, 16#06#),
      554 => to_slv(opcode_type, 16#09#),
      555 => to_slv(opcode_type, 16#0F#),
      556 => to_slv(opcode_type, 16#0F#),
      557 => to_slv(opcode_type, 16#06#),
      558 => to_slv(opcode_type, 16#0F#),
      559 => to_slv(opcode_type, 16#0B#),
      560 => to_slv(opcode_type, 16#09#),
      561 => to_slv(opcode_type, 16#08#),
      562 => to_slv(opcode_type, 16#09#),
      563 => to_slv(opcode_type, 16#11#),
      564 => to_slv(opcode_type, 16#0C#),
      565 => to_slv(opcode_type, 16#08#),
      566 => to_slv(opcode_type, 16#43#),
      567 => to_slv(opcode_type, 16#0A#),
      568 => to_slv(opcode_type, 16#08#),
      569 => to_slv(opcode_type, 16#08#),
      570 => to_slv(opcode_type, 16#BB#),
      571 => to_slv(opcode_type, 16#D7#),
      572 => to_slv(opcode_type, 16#08#),
      573 => to_slv(opcode_type, 16#0F#),
      574 => to_slv(opcode_type, 16#0F#),
      575 to 575 => (others => '0'),

      -- Program 18...
      576 => to_slv(opcode_type, 16#08#),
      577 => to_slv(opcode_type, 16#09#),
      578 => to_slv(opcode_type, 16#09#),
      579 => to_slv(opcode_type, 16#09#),
      580 => to_slv(opcode_type, 16#10#),
      581 => to_slv(opcode_type, 16#10#),
      582 => to_slv(opcode_type, 16#06#),
      583 => to_slv(opcode_type, 16#A4#),
      584 => to_slv(opcode_type, 16#0C#),
      585 => to_slv(opcode_type, 16#07#),
      586 => to_slv(opcode_type, 16#06#),
      587 => to_slv(opcode_type, 16#10#),
      588 => to_slv(opcode_type, 16#11#),
      589 => to_slv(opcode_type, 16#07#),
      590 => to_slv(opcode_type, 16#0F#),
      591 => to_slv(opcode_type, 16#0A#),
      592 => to_slv(opcode_type, 16#06#),
      593 => to_slv(opcode_type, 16#06#),
      594 => to_slv(opcode_type, 16#06#),
      595 => to_slv(opcode_type, 16#10#),
      596 => to_slv(opcode_type, 16#11#),
      597 => to_slv(opcode_type, 16#07#),
      598 => to_slv(opcode_type, 16#11#),
      599 => to_slv(opcode_type, 16#11#),
      600 => to_slv(opcode_type, 16#07#),
      601 => to_slv(opcode_type, 16#06#),
      602 => to_slv(opcode_type, 16#11#),
      603 => to_slv(opcode_type, 16#0D#),
      604 => to_slv(opcode_type, 16#09#),
      605 => to_slv(opcode_type, 16#11#),
      606 => to_slv(opcode_type, 16#83#),
      607 to 607 => (others => '0'),

      -- Program 19...
      608 => to_slv(opcode_type, 16#07#),
      609 => to_slv(opcode_type, 16#06#),
      610 => to_slv(opcode_type, 16#08#),
      611 => to_slv(opcode_type, 16#06#),
      612 => to_slv(opcode_type, 16#0B#),
      613 => to_slv(opcode_type, 16#11#),
      614 => to_slv(opcode_type, 16#09#),
      615 => to_slv(opcode_type, 16#0C#),
      616 => to_slv(opcode_type, 16#0B#),
      617 => to_slv(opcode_type, 16#09#),
      618 => to_slv(opcode_type, 16#08#),
      619 => to_slv(opcode_type, 16#0A#),
      620 => to_slv(opcode_type, 16#1C#),
      621 => to_slv(opcode_type, 16#09#),
      622 => to_slv(opcode_type, 16#0D#),
      623 => to_slv(opcode_type, 16#10#),
      624 => to_slv(opcode_type, 16#09#),
      625 => to_slv(opcode_type, 16#09#),
      626 => to_slv(opcode_type, 16#07#),
      627 => to_slv(opcode_type, 16#12#),
      628 => to_slv(opcode_type, 16#0F#),
      629 => to_slv(opcode_type, 16#08#),
      630 => to_slv(opcode_type, 16#11#),
      631 => to_slv(opcode_type, 16#0D#),
      632 => to_slv(opcode_type, 16#09#),
      633 => to_slv(opcode_type, 16#08#),
      634 => to_slv(opcode_type, 16#0B#),
      635 => to_slv(opcode_type, 16#0D#),
      636 => to_slv(opcode_type, 16#08#),
      637 => to_slv(opcode_type, 16#0F#),
      638 => to_slv(opcode_type, 16#D8#),
      639 to 639 => (others => '0'),

      -- Program 20...
      640 => to_slv(opcode_type, 16#09#),
      641 => to_slv(opcode_type, 16#07#),
      642 => to_slv(opcode_type, 16#09#),
      643 => to_slv(opcode_type, 16#06#),
      644 => to_slv(opcode_type, 16#AD#),
      645 => to_slv(opcode_type, 16#11#),
      646 => to_slv(opcode_type, 16#08#),
      647 => to_slv(opcode_type, 16#10#),
      648 => to_slv(opcode_type, 16#0C#),
      649 => to_slv(opcode_type, 16#06#),
      650 => to_slv(opcode_type, 16#07#),
      651 => to_slv(opcode_type, 16#11#),
      652 => to_slv(opcode_type, 16#10#),
      653 => to_slv(opcode_type, 16#06#),
      654 => to_slv(opcode_type, 16#11#),
      655 => to_slv(opcode_type, 16#37#),
      656 => to_slv(opcode_type, 16#08#),
      657 => to_slv(opcode_type, 16#06#),
      658 => to_slv(opcode_type, 16#06#),
      659 => to_slv(opcode_type, 16#0C#),
      660 => to_slv(opcode_type, 16#0E#),
      661 => to_slv(opcode_type, 16#06#),
      662 => to_slv(opcode_type, 16#11#),
      663 => to_slv(opcode_type, 16#0B#),
      664 => to_slv(opcode_type, 16#07#),
      665 => to_slv(opcode_type, 16#09#),
      666 => to_slv(opcode_type, 16#0E#),
      667 => to_slv(opcode_type, 16#0E#),
      668 => to_slv(opcode_type, 16#06#),
      669 => to_slv(opcode_type, 16#0A#),
      670 => to_slv(opcode_type, 16#10#),
      671 to 671 => (others => '0'),

      -- Program 21...
      672 => to_slv(opcode_type, 16#07#),
      673 => to_slv(opcode_type, 16#08#),
      674 => to_slv(opcode_type, 16#09#),
      675 => to_slv(opcode_type, 16#06#),
      676 => to_slv(opcode_type, 16#10#),
      677 => to_slv(opcode_type, 16#0D#),
      678 => to_slv(opcode_type, 16#08#),
      679 => to_slv(opcode_type, 16#0A#),
      680 => to_slv(opcode_type, 16#91#),
      681 => to_slv(opcode_type, 16#08#),
      682 => to_slv(opcode_type, 16#07#),
      683 => to_slv(opcode_type, 16#10#),
      684 => to_slv(opcode_type, 16#0B#),
      685 => to_slv(opcode_type, 16#07#),
      686 => to_slv(opcode_type, 16#0A#),
      687 => to_slv(opcode_type, 16#10#),
      688 => to_slv(opcode_type, 16#09#),
      689 => to_slv(opcode_type, 16#08#),
      690 => to_slv(opcode_type, 16#06#),
      691 => to_slv(opcode_type, 16#0D#),
      692 => to_slv(opcode_type, 16#0F#),
      693 => to_slv(opcode_type, 16#09#),
      694 => to_slv(opcode_type, 16#0A#),
      695 => to_slv(opcode_type, 16#0E#),
      696 => to_slv(opcode_type, 16#09#),
      697 => to_slv(opcode_type, 16#06#),
      698 => to_slv(opcode_type, 16#0E#),
      699 => to_slv(opcode_type, 16#0F#),
      700 => to_slv(opcode_type, 16#07#),
      701 => to_slv(opcode_type, 16#11#),
      702 => to_slv(opcode_type, 16#11#),
      703 to 703 => (others => '0'),

      -- Program 22...
      704 => to_slv(opcode_type, 16#09#),
      705 => to_slv(opcode_type, 16#08#),
      706 => to_slv(opcode_type, 16#09#),
      707 => to_slv(opcode_type, 16#07#),
      708 => to_slv(opcode_type, 16#0B#),
      709 => to_slv(opcode_type, 16#0E#),
      710 => to_slv(opcode_type, 16#06#),
      711 => to_slv(opcode_type, 16#0F#),
      712 => to_slv(opcode_type, 16#0C#),
      713 => to_slv(opcode_type, 16#09#),
      714 => to_slv(opcode_type, 16#08#),
      715 => to_slv(opcode_type, 16#0B#),
      716 => to_slv(opcode_type, 16#0E#),
      717 => to_slv(opcode_type, 16#07#),
      718 => to_slv(opcode_type, 16#0E#),
      719 => to_slv(opcode_type, 16#10#),
      720 => to_slv(opcode_type, 16#07#),
      721 => to_slv(opcode_type, 16#09#),
      722 => to_slv(opcode_type, 16#07#),
      723 => to_slv(opcode_type, 16#0B#),
      724 => to_slv(opcode_type, 16#10#),
      725 => to_slv(opcode_type, 16#07#),
      726 => to_slv(opcode_type, 16#0B#),
      727 => to_slv(opcode_type, 16#0C#),
      728 => to_slv(opcode_type, 16#08#),
      729 => to_slv(opcode_type, 16#07#),
      730 => to_slv(opcode_type, 16#0C#),
      731 => to_slv(opcode_type, 16#0F#),
      732 => to_slv(opcode_type, 16#07#),
      733 => to_slv(opcode_type, 16#0F#),
      734 => to_slv(opcode_type, 16#0E#),
      735 to 735 => (others => '0'),

      -- Program 23...
      736 => to_slv(opcode_type, 16#09#),
      737 => to_slv(opcode_type, 16#06#),
      738 => to_slv(opcode_type, 16#07#),
      739 => to_slv(opcode_type, 16#08#),
      740 => to_slv(opcode_type, 16#0F#),
      741 => to_slv(opcode_type, 16#0D#),
      742 => to_slv(opcode_type, 16#08#),
      743 => to_slv(opcode_type, 16#0C#),
      744 => to_slv(opcode_type, 16#11#),
      745 => to_slv(opcode_type, 16#07#),
      746 => to_slv(opcode_type, 16#08#),
      747 => to_slv(opcode_type, 16#0F#),
      748 => to_slv(opcode_type, 16#11#),
      749 => to_slv(opcode_type, 16#06#),
      750 => to_slv(opcode_type, 16#0B#),
      751 => to_slv(opcode_type, 16#0D#),
      752 => to_slv(opcode_type, 16#06#),
      753 => to_slv(opcode_type, 16#06#),
      754 => to_slv(opcode_type, 16#06#),
      755 => to_slv(opcode_type, 16#0E#),
      756 => to_slv(opcode_type, 16#10#),
      757 => to_slv(opcode_type, 16#08#),
      758 => to_slv(opcode_type, 16#0A#),
      759 => to_slv(opcode_type, 16#0A#),
      760 => to_slv(opcode_type, 16#09#),
      761 => to_slv(opcode_type, 16#07#),
      762 => to_slv(opcode_type, 16#0B#),
      763 => to_slv(opcode_type, 16#0E#),
      764 => to_slv(opcode_type, 16#08#),
      765 => to_slv(opcode_type, 16#DD#),
      766 => to_slv(opcode_type, 16#0C#),
      767 to 767 => (others => '0'),

      -- Program 24...
      768 => to_slv(opcode_type, 16#08#),
      769 => to_slv(opcode_type, 16#08#),
      770 => to_slv(opcode_type, 16#07#),
      771 => to_slv(opcode_type, 16#06#),
      772 => to_slv(opcode_type, 16#0B#),
      773 => to_slv(opcode_type, 16#10#),
      774 => to_slv(opcode_type, 16#08#),
      775 => to_slv(opcode_type, 16#0A#),
      776 => to_slv(opcode_type, 16#0E#),
      777 => to_slv(opcode_type, 16#09#),
      778 => to_slv(opcode_type, 16#08#),
      779 => to_slv(opcode_type, 16#C7#),
      780 => to_slv(opcode_type, 16#C1#),
      781 => to_slv(opcode_type, 16#09#),
      782 => to_slv(opcode_type, 16#0D#),
      783 => to_slv(opcode_type, 16#10#),
      784 => to_slv(opcode_type, 16#06#),
      785 => to_slv(opcode_type, 16#08#),
      786 => to_slv(opcode_type, 16#06#),
      787 => to_slv(opcode_type, 16#10#),
      788 => to_slv(opcode_type, 16#0F#),
      789 => to_slv(opcode_type, 16#07#),
      790 => to_slv(opcode_type, 16#0D#),
      791 => to_slv(opcode_type, 16#0B#),
      792 => to_slv(opcode_type, 16#07#),
      793 => to_slv(opcode_type, 16#08#),
      794 => to_slv(opcode_type, 16#0B#),
      795 => to_slv(opcode_type, 16#0E#),
      796 => to_slv(opcode_type, 16#06#),
      797 => to_slv(opcode_type, 16#0D#),
      798 => to_slv(opcode_type, 16#0B#),
      799 to 799 => (others => '0'),

      -- Program 25...
      800 => to_slv(opcode_type, 16#08#),
      801 => to_slv(opcode_type, 16#08#),
      802 => to_slv(opcode_type, 16#07#),
      803 => to_slv(opcode_type, 16#06#),
      804 => to_slv(opcode_type, 16#AD#),
      805 => to_slv(opcode_type, 16#0D#),
      806 => to_slv(opcode_type, 16#09#),
      807 => to_slv(opcode_type, 16#0D#),
      808 => to_slv(opcode_type, 16#0A#),
      809 => to_slv(opcode_type, 16#08#),
      810 => to_slv(opcode_type, 16#09#),
      811 => to_slv(opcode_type, 16#0A#),
      812 => to_slv(opcode_type, 16#0B#),
      813 => to_slv(opcode_type, 16#07#),
      814 => to_slv(opcode_type, 16#0F#),
      815 => to_slv(opcode_type, 16#0F#),
      816 => to_slv(opcode_type, 16#08#),
      817 => to_slv(opcode_type, 16#06#),
      818 => to_slv(opcode_type, 16#08#),
      819 => to_slv(opcode_type, 16#10#),
      820 => to_slv(opcode_type, 16#0D#),
      821 => to_slv(opcode_type, 16#08#),
      822 => to_slv(opcode_type, 16#0B#),
      823 => to_slv(opcode_type, 16#11#),
      824 => to_slv(opcode_type, 16#08#),
      825 => to_slv(opcode_type, 16#07#),
      826 => to_slv(opcode_type, 16#0E#),
      827 => to_slv(opcode_type, 16#11#),
      828 => to_slv(opcode_type, 16#09#),
      829 => to_slv(opcode_type, 16#0E#),
      830 => to_slv(opcode_type, 16#11#),
      831 to 831 => (others => '0'),

      -- Program 26...
      832 => to_slv(opcode_type, 16#07#),
      833 => to_slv(opcode_type, 16#07#),
      834 => to_slv(opcode_type, 16#08#),
      835 => to_slv(opcode_type, 16#09#),
      836 => to_slv(opcode_type, 16#0C#),
      837 => to_slv(opcode_type, 16#0B#),
      838 => to_slv(opcode_type, 16#09#),
      839 => to_slv(opcode_type, 16#0C#),
      840 => to_slv(opcode_type, 16#0F#),
      841 => to_slv(opcode_type, 16#09#),
      842 => to_slv(opcode_type, 16#08#),
      843 => to_slv(opcode_type, 16#0C#),
      844 => to_slv(opcode_type, 16#A3#),
      845 => to_slv(opcode_type, 16#07#),
      846 => to_slv(opcode_type, 16#54#),
      847 => to_slv(opcode_type, 16#0C#),
      848 => to_slv(opcode_type, 16#07#),
      849 => to_slv(opcode_type, 16#06#),
      850 => to_slv(opcode_type, 16#07#),
      851 => to_slv(opcode_type, 16#0A#),
      852 => to_slv(opcode_type, 16#0D#),
      853 => to_slv(opcode_type, 16#09#),
      854 => to_slv(opcode_type, 16#0B#),
      855 => to_slv(opcode_type, 16#0F#),
      856 => to_slv(opcode_type, 16#06#),
      857 => to_slv(opcode_type, 16#09#),
      858 => to_slv(opcode_type, 16#11#),
      859 => to_slv(opcode_type, 16#0A#),
      860 => to_slv(opcode_type, 16#09#),
      861 => to_slv(opcode_type, 16#0F#),
      862 => to_slv(opcode_type, 16#0D#),
      863 to 863 => (others => '0'),

      -- Program 27...
      864 => to_slv(opcode_type, 16#09#),
      865 => to_slv(opcode_type, 16#09#),
      866 => to_slv(opcode_type, 16#09#),
      867 => to_slv(opcode_type, 16#08#),
      868 => to_slv(opcode_type, 16#0C#),
      869 => to_slv(opcode_type, 16#0D#),
      870 => to_slv(opcode_type, 16#09#),
      871 => to_slv(opcode_type, 16#0D#),
      872 => to_slv(opcode_type, 16#0C#),
      873 => to_slv(opcode_type, 16#07#),
      874 => to_slv(opcode_type, 16#07#),
      875 => to_slv(opcode_type, 16#0A#),
      876 => to_slv(opcode_type, 16#11#),
      877 => to_slv(opcode_type, 16#07#),
      878 => to_slv(opcode_type, 16#11#),
      879 => to_slv(opcode_type, 16#0F#),
      880 => to_slv(opcode_type, 16#06#),
      881 => to_slv(opcode_type, 16#07#),
      882 => to_slv(opcode_type, 16#06#),
      883 => to_slv(opcode_type, 16#0F#),
      884 => to_slv(opcode_type, 16#11#),
      885 => to_slv(opcode_type, 16#08#),
      886 => to_slv(opcode_type, 16#11#),
      887 => to_slv(opcode_type, 16#C6#),
      888 => to_slv(opcode_type, 16#06#),
      889 => to_slv(opcode_type, 16#08#),
      890 => to_slv(opcode_type, 16#10#),
      891 => to_slv(opcode_type, 16#0A#),
      892 => to_slv(opcode_type, 16#06#),
      893 => to_slv(opcode_type, 16#0D#),
      894 => to_slv(opcode_type, 16#70#),
      895 to 895 => (others => '0'),

      -- Program 28...
      896 => to_slv(opcode_type, 16#06#),
      897 => to_slv(opcode_type, 16#08#),
      898 => to_slv(opcode_type, 16#06#),
      899 => to_slv(opcode_type, 16#08#),
      900 => to_slv(opcode_type, 16#0A#),
      901 => to_slv(opcode_type, 16#0D#),
      902 => to_slv(opcode_type, 16#07#),
      903 => to_slv(opcode_type, 16#0A#),
      904 => to_slv(opcode_type, 16#0F#),
      905 => to_slv(opcode_type, 16#07#),
      906 => to_slv(opcode_type, 16#06#),
      907 => to_slv(opcode_type, 16#0A#),
      908 => to_slv(opcode_type, 16#10#),
      909 => to_slv(opcode_type, 16#08#),
      910 => to_slv(opcode_type, 16#0A#),
      911 => to_slv(opcode_type, 16#0A#),
      912 => to_slv(opcode_type, 16#06#),
      913 => to_slv(opcode_type, 16#07#),
      914 => to_slv(opcode_type, 16#09#),
      915 => to_slv(opcode_type, 16#0F#),
      916 => to_slv(opcode_type, 16#11#),
      917 => to_slv(opcode_type, 16#09#),
      918 => to_slv(opcode_type, 16#B5#),
      919 => to_slv(opcode_type, 16#0B#),
      920 => to_slv(opcode_type, 16#08#),
      921 => to_slv(opcode_type, 16#07#),
      922 => to_slv(opcode_type, 16#10#),
      923 => to_slv(opcode_type, 16#10#),
      924 => to_slv(opcode_type, 16#07#),
      925 => to_slv(opcode_type, 16#0D#),
      926 => to_slv(opcode_type, 16#0E#),
      927 to 927 => (others => '0'),

      -- Program 29...
      928 => to_slv(opcode_type, 16#09#),
      929 => to_slv(opcode_type, 16#09#),
      930 => to_slv(opcode_type, 16#08#),
      931 => to_slv(opcode_type, 16#07#),
      932 => to_slv(opcode_type, 16#0C#),
      933 => to_slv(opcode_type, 16#0A#),
      934 => to_slv(opcode_type, 16#09#),
      935 => to_slv(opcode_type, 16#9E#),
      936 => to_slv(opcode_type, 16#10#),
      937 => to_slv(opcode_type, 16#08#),
      938 => to_slv(opcode_type, 16#07#),
      939 => to_slv(opcode_type, 16#0F#),
      940 => to_slv(opcode_type, 16#0E#),
      941 => to_slv(opcode_type, 16#07#),
      942 => to_slv(opcode_type, 16#0E#),
      943 => to_slv(opcode_type, 16#11#),
      944 => to_slv(opcode_type, 16#07#),
      945 => to_slv(opcode_type, 16#08#),
      946 => to_slv(opcode_type, 16#07#),
      947 => to_slv(opcode_type, 16#0D#),
      948 => to_slv(opcode_type, 16#0D#),
      949 => to_slv(opcode_type, 16#08#),
      950 => to_slv(opcode_type, 16#20#),
      951 => to_slv(opcode_type, 16#0B#),
      952 => to_slv(opcode_type, 16#08#),
      953 => to_slv(opcode_type, 16#06#),
      954 => to_slv(opcode_type, 16#0B#),
      955 => to_slv(opcode_type, 16#10#),
      956 => to_slv(opcode_type, 16#08#),
      957 => to_slv(opcode_type, 16#0A#),
      958 => to_slv(opcode_type, 16#0A#),
      959 to 959 => (others => '0'),

      -- Program 30...
      960 => to_slv(opcode_type, 16#08#),
      961 => to_slv(opcode_type, 16#06#),
      962 => to_slv(opcode_type, 16#07#),
      963 => to_slv(opcode_type, 16#09#),
      964 => to_slv(opcode_type, 16#46#),
      965 => to_slv(opcode_type, 16#0B#),
      966 => to_slv(opcode_type, 16#06#),
      967 => to_slv(opcode_type, 16#0B#),
      968 => to_slv(opcode_type, 16#0D#),
      969 => to_slv(opcode_type, 16#08#),
      970 => to_slv(opcode_type, 16#07#),
      971 => to_slv(opcode_type, 16#1F#),
      972 => to_slv(opcode_type, 16#BD#),
      973 => to_slv(opcode_type, 16#07#),
      974 => to_slv(opcode_type, 16#11#),
      975 => to_slv(opcode_type, 16#0C#),
      976 => to_slv(opcode_type, 16#08#),
      977 => to_slv(opcode_type, 16#07#),
      978 => to_slv(opcode_type, 16#09#),
      979 => to_slv(opcode_type, 16#11#),
      980 => to_slv(opcode_type, 16#0B#),
      981 => to_slv(opcode_type, 16#09#),
      982 => to_slv(opcode_type, 16#0A#),
      983 => to_slv(opcode_type, 16#0A#),
      984 => to_slv(opcode_type, 16#07#),
      985 => to_slv(opcode_type, 16#06#),
      986 => to_slv(opcode_type, 16#0D#),
      987 => to_slv(opcode_type, 16#0C#),
      988 => to_slv(opcode_type, 16#06#),
      989 => to_slv(opcode_type, 16#BC#),
      990 => to_slv(opcode_type, 16#11#),
      991 to 991 => (others => '0'),

      -- Program 31...
      992 => to_slv(opcode_type, 16#08#),
      993 => to_slv(opcode_type, 16#09#),
      994 => to_slv(opcode_type, 16#09#),
      995 => to_slv(opcode_type, 16#08#),
      996 => to_slv(opcode_type, 16#45#),
      997 => to_slv(opcode_type, 16#0A#),
      998 => to_slv(opcode_type, 16#08#),
      999 => to_slv(opcode_type, 16#0B#),
      1000 => to_slv(opcode_type, 16#10#),
      1001 => to_slv(opcode_type, 16#09#),
      1002 => to_slv(opcode_type, 16#09#),
      1003 => to_slv(opcode_type, 16#0D#),
      1004 => to_slv(opcode_type, 16#11#),
      1005 => to_slv(opcode_type, 16#07#),
      1006 => to_slv(opcode_type, 16#10#),
      1007 => to_slv(opcode_type, 16#10#),
      1008 => to_slv(opcode_type, 16#07#),
      1009 => to_slv(opcode_type, 16#07#),
      1010 => to_slv(opcode_type, 16#07#),
      1011 => to_slv(opcode_type, 16#0B#),
      1012 => to_slv(opcode_type, 16#0D#),
      1013 => to_slv(opcode_type, 16#06#),
      1014 => to_slv(opcode_type, 16#10#),
      1015 => to_slv(opcode_type, 16#0F#),
      1016 => to_slv(opcode_type, 16#09#),
      1017 => to_slv(opcode_type, 16#08#),
      1018 => to_slv(opcode_type, 16#0A#),
      1019 => to_slv(opcode_type, 16#11#),
      1020 => to_slv(opcode_type, 16#08#),
      1021 => to_slv(opcode_type, 16#0D#),
      1022 => to_slv(opcode_type, 16#0A#),
      1023 to 1023 => (others => '0'),

      -- Program 32...
      1024 => to_slv(opcode_type, 16#06#),
      1025 => to_slv(opcode_type, 16#08#),
      1026 => to_slv(opcode_type, 16#07#),
      1027 => to_slv(opcode_type, 16#07#),
      1028 => to_slv(opcode_type, 16#0B#),
      1029 => to_slv(opcode_type, 16#0E#),
      1030 => to_slv(opcode_type, 16#07#),
      1031 => to_slv(opcode_type, 16#0D#),
      1032 => to_slv(opcode_type, 16#0B#),
      1033 => to_slv(opcode_type, 16#07#),
      1034 => to_slv(opcode_type, 16#08#),
      1035 => to_slv(opcode_type, 16#0D#),
      1036 => to_slv(opcode_type, 16#10#),
      1037 => to_slv(opcode_type, 16#09#),
      1038 => to_slv(opcode_type, 16#0C#),
      1039 => to_slv(opcode_type, 16#0A#),
      1040 => to_slv(opcode_type, 16#07#),
      1041 => to_slv(opcode_type, 16#06#),
      1042 => to_slv(opcode_type, 16#08#),
      1043 => to_slv(opcode_type, 16#1F#),
      1044 => to_slv(opcode_type, 16#0D#),
      1045 => to_slv(opcode_type, 16#07#),
      1046 => to_slv(opcode_type, 16#11#),
      1047 => to_slv(opcode_type, 16#0F#),
      1048 => to_slv(opcode_type, 16#09#),
      1049 => to_slv(opcode_type, 16#06#),
      1050 => to_slv(opcode_type, 16#0C#),
      1051 => to_slv(opcode_type, 16#10#),
      1052 => to_slv(opcode_type, 16#09#),
      1053 => to_slv(opcode_type, 16#0E#),
      1054 => to_slv(opcode_type, 16#0C#),
      1055 to 1055 => (others => '0'),

      -- Program 33...
      1056 => to_slv(opcode_type, 16#06#),
      1057 => to_slv(opcode_type, 16#07#),
      1058 => to_slv(opcode_type, 16#08#),
      1059 => to_slv(opcode_type, 16#06#),
      1060 => to_slv(opcode_type, 16#11#),
      1061 => to_slv(opcode_type, 16#0D#),
      1062 => to_slv(opcode_type, 16#06#),
      1063 => to_slv(opcode_type, 16#0A#),
      1064 => to_slv(opcode_type, 16#0D#),
      1065 => to_slv(opcode_type, 16#08#),
      1066 => to_slv(opcode_type, 16#06#),
      1067 => to_slv(opcode_type, 16#0C#),
      1068 => to_slv(opcode_type, 16#0E#),
      1069 => to_slv(opcode_type, 16#07#),
      1070 => to_slv(opcode_type, 16#D8#),
      1071 => to_slv(opcode_type, 16#0C#),
      1072 => to_slv(opcode_type, 16#08#),
      1073 => to_slv(opcode_type, 16#08#),
      1074 => to_slv(opcode_type, 16#06#),
      1075 => to_slv(opcode_type, 16#0E#),
      1076 => to_slv(opcode_type, 16#0A#),
      1077 => to_slv(opcode_type, 16#07#),
      1078 => to_slv(opcode_type, 16#0E#),
      1079 => to_slv(opcode_type, 16#0B#),
      1080 => to_slv(opcode_type, 16#09#),
      1081 => to_slv(opcode_type, 16#08#),
      1082 => to_slv(opcode_type, 16#0F#),
      1083 => to_slv(opcode_type, 16#0F#),
      1084 => to_slv(opcode_type, 16#07#),
      1085 => to_slv(opcode_type, 16#11#),
      1086 => to_slv(opcode_type, 16#0C#),
      1087 to 1087 => (others => '0'),

      -- Program 34...
      1088 => to_slv(opcode_type, 16#06#),
      1089 => to_slv(opcode_type, 16#07#),
      1090 => to_slv(opcode_type, 16#07#),
      1091 => to_slv(opcode_type, 16#06#),
      1092 => to_slv(opcode_type, 16#0D#),
      1093 => to_slv(opcode_type, 16#10#),
      1094 => to_slv(opcode_type, 16#08#),
      1095 => to_slv(opcode_type, 16#0F#),
      1096 => to_slv(opcode_type, 16#0D#),
      1097 => to_slv(opcode_type, 16#07#),
      1098 => to_slv(opcode_type, 16#08#),
      1099 => to_slv(opcode_type, 16#0A#),
      1100 => to_slv(opcode_type, 16#0E#),
      1101 => to_slv(opcode_type, 16#07#),
      1102 => to_slv(opcode_type, 16#0B#),
      1103 => to_slv(opcode_type, 16#0D#),
      1104 => to_slv(opcode_type, 16#09#),
      1105 => to_slv(opcode_type, 16#08#),
      1106 => to_slv(opcode_type, 16#06#),
      1107 => to_slv(opcode_type, 16#0E#),
      1108 => to_slv(opcode_type, 16#0E#),
      1109 => to_slv(opcode_type, 16#06#),
      1110 => to_slv(opcode_type, 16#0F#),
      1111 => to_slv(opcode_type, 16#8E#),
      1112 => to_slv(opcode_type, 16#06#),
      1113 => to_slv(opcode_type, 16#07#),
      1114 => to_slv(opcode_type, 16#0D#),
      1115 => to_slv(opcode_type, 16#0A#),
      1116 => to_slv(opcode_type, 16#07#),
      1117 => to_slv(opcode_type, 16#0D#),
      1118 => to_slv(opcode_type, 16#0C#),
      1119 to 1119 => (others => '0'),

      -- Program 35...
      1120 => to_slv(opcode_type, 16#07#),
      1121 => to_slv(opcode_type, 16#09#),
      1122 => to_slv(opcode_type, 16#08#),
      1123 => to_slv(opcode_type, 16#08#),
      1124 => to_slv(opcode_type, 16#10#),
      1125 => to_slv(opcode_type, 16#0D#),
      1126 => to_slv(opcode_type, 16#07#),
      1127 => to_slv(opcode_type, 16#10#),
      1128 => to_slv(opcode_type, 16#0E#),
      1129 => to_slv(opcode_type, 16#08#),
      1130 => to_slv(opcode_type, 16#06#),
      1131 => to_slv(opcode_type, 16#10#),
      1132 => to_slv(opcode_type, 16#0D#),
      1133 => to_slv(opcode_type, 16#08#),
      1134 => to_slv(opcode_type, 16#0E#),
      1135 => to_slv(opcode_type, 16#0C#),
      1136 => to_slv(opcode_type, 16#07#),
      1137 => to_slv(opcode_type, 16#08#),
      1138 => to_slv(opcode_type, 16#06#),
      1139 => to_slv(opcode_type, 16#0C#),
      1140 => to_slv(opcode_type, 16#10#),
      1141 => to_slv(opcode_type, 16#08#),
      1142 => to_slv(opcode_type, 16#11#),
      1143 => to_slv(opcode_type, 16#0C#),
      1144 => to_slv(opcode_type, 16#07#),
      1145 => to_slv(opcode_type, 16#09#),
      1146 => to_slv(opcode_type, 16#0F#),
      1147 => to_slv(opcode_type, 16#10#),
      1148 => to_slv(opcode_type, 16#06#),
      1149 => to_slv(opcode_type, 16#0A#),
      1150 => to_slv(opcode_type, 16#0B#),
      1151 to 1151 => (others => '0'),

      -- Program 36...
      1152 => to_slv(opcode_type, 16#06#),
      1153 => to_slv(opcode_type, 16#09#),
      1154 => to_slv(opcode_type, 16#08#),
      1155 => to_slv(opcode_type, 16#08#),
      1156 => to_slv(opcode_type, 16#0C#),
      1157 => to_slv(opcode_type, 16#0A#),
      1158 => to_slv(opcode_type, 16#06#),
      1159 => to_slv(opcode_type, 16#0A#),
      1160 => to_slv(opcode_type, 16#0E#),
      1161 => to_slv(opcode_type, 16#09#),
      1162 => to_slv(opcode_type, 16#09#),
      1163 => to_slv(opcode_type, 16#0C#),
      1164 => to_slv(opcode_type, 16#0C#),
      1165 => to_slv(opcode_type, 16#09#),
      1166 => to_slv(opcode_type, 16#0E#),
      1167 => to_slv(opcode_type, 16#0E#),
      1168 => to_slv(opcode_type, 16#09#),
      1169 => to_slv(opcode_type, 16#07#),
      1170 => to_slv(opcode_type, 16#09#),
      1171 => to_slv(opcode_type, 16#0E#),
      1172 => to_slv(opcode_type, 16#0A#),
      1173 => to_slv(opcode_type, 16#08#),
      1174 => to_slv(opcode_type, 16#10#),
      1175 => to_slv(opcode_type, 16#0D#),
      1176 => to_slv(opcode_type, 16#07#),
      1177 => to_slv(opcode_type, 16#08#),
      1178 => to_slv(opcode_type, 16#0C#),
      1179 => to_slv(opcode_type, 16#10#),
      1180 => to_slv(opcode_type, 16#06#),
      1181 => to_slv(opcode_type, 16#10#),
      1182 => to_slv(opcode_type, 16#0C#),
      1183 to 1183 => (others => '0'),

      -- Program 37...
      1184 => to_slv(opcode_type, 16#06#),
      1185 => to_slv(opcode_type, 16#07#),
      1186 => to_slv(opcode_type, 16#07#),
      1187 => to_slv(opcode_type, 16#08#),
      1188 => to_slv(opcode_type, 16#0C#),
      1189 => to_slv(opcode_type, 16#54#),
      1190 => to_slv(opcode_type, 16#09#),
      1191 => to_slv(opcode_type, 16#0D#),
      1192 => to_slv(opcode_type, 16#0D#),
      1193 => to_slv(opcode_type, 16#07#),
      1194 => to_slv(opcode_type, 16#09#),
      1195 => to_slv(opcode_type, 16#0A#),
      1196 => to_slv(opcode_type, 16#0F#),
      1197 => to_slv(opcode_type, 16#09#),
      1198 => to_slv(opcode_type, 16#0B#),
      1199 => to_slv(opcode_type, 16#0F#),
      1200 => to_slv(opcode_type, 16#07#),
      1201 => to_slv(opcode_type, 16#06#),
      1202 => to_slv(opcode_type, 16#07#),
      1203 => to_slv(opcode_type, 16#0E#),
      1204 => to_slv(opcode_type, 16#0F#),
      1205 => to_slv(opcode_type, 16#07#),
      1206 => to_slv(opcode_type, 16#0F#),
      1207 => to_slv(opcode_type, 16#0F#),
      1208 => to_slv(opcode_type, 16#08#),
      1209 => to_slv(opcode_type, 16#09#),
      1210 => to_slv(opcode_type, 16#0A#),
      1211 => to_slv(opcode_type, 16#0A#),
      1212 => to_slv(opcode_type, 16#06#),
      1213 => to_slv(opcode_type, 16#11#),
      1214 => to_slv(opcode_type, 16#0A#),
      1215 to 1215 => (others => '0'),

      -- Program 38...
      1216 => to_slv(opcode_type, 16#06#),
      1217 => to_slv(opcode_type, 16#09#),
      1218 => to_slv(opcode_type, 16#07#),
      1219 => to_slv(opcode_type, 16#09#),
      1220 => to_slv(opcode_type, 16#0D#),
      1221 => to_slv(opcode_type, 16#0F#),
      1222 => to_slv(opcode_type, 16#08#),
      1223 => to_slv(opcode_type, 16#2A#),
      1224 => to_slv(opcode_type, 16#0E#),
      1225 => to_slv(opcode_type, 16#09#),
      1226 => to_slv(opcode_type, 16#06#),
      1227 => to_slv(opcode_type, 16#0B#),
      1228 => to_slv(opcode_type, 16#10#),
      1229 => to_slv(opcode_type, 16#06#),
      1230 => to_slv(opcode_type, 16#0F#),
      1231 => to_slv(opcode_type, 16#0C#),
      1232 => to_slv(opcode_type, 16#09#),
      1233 => to_slv(opcode_type, 16#06#),
      1234 => to_slv(opcode_type, 16#06#),
      1235 => to_slv(opcode_type, 16#0F#),
      1236 => to_slv(opcode_type, 16#0B#),
      1237 => to_slv(opcode_type, 16#06#),
      1238 => to_slv(opcode_type, 16#10#),
      1239 => to_slv(opcode_type, 16#10#),
      1240 => to_slv(opcode_type, 16#07#),
      1241 => to_slv(opcode_type, 16#07#),
      1242 => to_slv(opcode_type, 16#0D#),
      1243 => to_slv(opcode_type, 16#C0#),
      1244 => to_slv(opcode_type, 16#08#),
      1245 => to_slv(opcode_type, 16#E9#),
      1246 => to_slv(opcode_type, 16#0B#),
      1247 to 1247 => (others => '0'),

      -- Program 39...
      1248 => to_slv(opcode_type, 16#08#),
      1249 => to_slv(opcode_type, 16#06#),
      1250 => to_slv(opcode_type, 16#06#),
      1251 => to_slv(opcode_type, 16#09#),
      1252 => to_slv(opcode_type, 16#0C#),
      1253 => to_slv(opcode_type, 16#0E#),
      1254 => to_slv(opcode_type, 16#09#),
      1255 => to_slv(opcode_type, 16#0B#),
      1256 => to_slv(opcode_type, 16#E0#),
      1257 => to_slv(opcode_type, 16#08#),
      1258 => to_slv(opcode_type, 16#09#),
      1259 => to_slv(opcode_type, 16#11#),
      1260 => to_slv(opcode_type, 16#0B#),
      1261 => to_slv(opcode_type, 16#07#),
      1262 => to_slv(opcode_type, 16#0E#),
      1263 => to_slv(opcode_type, 16#10#),
      1264 => to_slv(opcode_type, 16#06#),
      1265 => to_slv(opcode_type, 16#06#),
      1266 => to_slv(opcode_type, 16#08#),
      1267 => to_slv(opcode_type, 16#0B#),
      1268 => to_slv(opcode_type, 16#0E#),
      1269 => to_slv(opcode_type, 16#08#),
      1270 => to_slv(opcode_type, 16#0F#),
      1271 => to_slv(opcode_type, 16#F7#),
      1272 => to_slv(opcode_type, 16#09#),
      1273 => to_slv(opcode_type, 16#08#),
      1274 => to_slv(opcode_type, 16#0A#),
      1275 => to_slv(opcode_type, 16#0E#),
      1276 => to_slv(opcode_type, 16#07#),
      1277 => to_slv(opcode_type, 16#0F#),
      1278 => to_slv(opcode_type, 16#0C#),
      1279 to 1279 => (others => '0'),

      -- Program 40...
      1280 => to_slv(opcode_type, 16#06#),
      1281 => to_slv(opcode_type, 16#07#),
      1282 => to_slv(opcode_type, 16#07#),
      1283 => to_slv(opcode_type, 16#08#),
      1284 => to_slv(opcode_type, 16#11#),
      1285 => to_slv(opcode_type, 16#13#),
      1286 => to_slv(opcode_type, 16#07#),
      1287 => to_slv(opcode_type, 16#11#),
      1288 => to_slv(opcode_type, 16#0D#),
      1289 => to_slv(opcode_type, 16#06#),
      1290 => to_slv(opcode_type, 16#07#),
      1291 => to_slv(opcode_type, 16#0F#),
      1292 => to_slv(opcode_type, 16#0C#),
      1293 => to_slv(opcode_type, 16#08#),
      1294 => to_slv(opcode_type, 16#10#),
      1295 => to_slv(opcode_type, 16#0B#),
      1296 => to_slv(opcode_type, 16#09#),
      1297 => to_slv(opcode_type, 16#09#),
      1298 => to_slv(opcode_type, 16#06#),
      1299 => to_slv(opcode_type, 16#10#),
      1300 => to_slv(opcode_type, 16#0D#),
      1301 => to_slv(opcode_type, 16#06#),
      1302 => to_slv(opcode_type, 16#A5#),
      1303 => to_slv(opcode_type, 16#0D#),
      1304 => to_slv(opcode_type, 16#09#),
      1305 => to_slv(opcode_type, 16#07#),
      1306 => to_slv(opcode_type, 16#D7#),
      1307 => to_slv(opcode_type, 16#10#),
      1308 => to_slv(opcode_type, 16#06#),
      1309 => to_slv(opcode_type, 16#44#),
      1310 => to_slv(opcode_type, 16#0F#),
      1311 to 1311 => (others => '0'),

      -- Program 41...
      1312 => to_slv(opcode_type, 16#06#),
      1313 => to_slv(opcode_type, 16#06#),
      1314 => to_slv(opcode_type, 16#06#),
      1315 => to_slv(opcode_type, 16#06#),
      1316 => to_slv(opcode_type, 16#0C#),
      1317 => to_slv(opcode_type, 16#0A#),
      1318 => to_slv(opcode_type, 16#09#),
      1319 => to_slv(opcode_type, 16#11#),
      1320 => to_slv(opcode_type, 16#0B#),
      1321 => to_slv(opcode_type, 16#06#),
      1322 => to_slv(opcode_type, 16#06#),
      1323 => to_slv(opcode_type, 16#10#),
      1324 => to_slv(opcode_type, 16#0F#),
      1325 => to_slv(opcode_type, 16#08#),
      1326 => to_slv(opcode_type, 16#0A#),
      1327 => to_slv(opcode_type, 16#0F#),
      1328 => to_slv(opcode_type, 16#08#),
      1329 => to_slv(opcode_type, 16#09#),
      1330 => to_slv(opcode_type, 16#08#),
      1331 => to_slv(opcode_type, 16#0F#),
      1332 => to_slv(opcode_type, 16#11#),
      1333 => to_slv(opcode_type, 16#06#),
      1334 => to_slv(opcode_type, 16#0C#),
      1335 => to_slv(opcode_type, 16#0D#),
      1336 => to_slv(opcode_type, 16#06#),
      1337 => to_slv(opcode_type, 16#06#),
      1338 => to_slv(opcode_type, 16#0E#),
      1339 => to_slv(opcode_type, 16#0D#),
      1340 => to_slv(opcode_type, 16#09#),
      1341 => to_slv(opcode_type, 16#0F#),
      1342 => to_slv(opcode_type, 16#0C#),
      1343 to 1343 => (others => '0'),

      -- Program 42...
      1344 => to_slv(opcode_type, 16#07#),
      1345 => to_slv(opcode_type, 16#08#),
      1346 => to_slv(opcode_type, 16#08#),
      1347 => to_slv(opcode_type, 16#07#),
      1348 => to_slv(opcode_type, 16#0F#),
      1349 => to_slv(opcode_type, 16#0F#),
      1350 => to_slv(opcode_type, 16#09#),
      1351 => to_slv(opcode_type, 16#F8#),
      1352 => to_slv(opcode_type, 16#0C#),
      1353 => to_slv(opcode_type, 16#09#),
      1354 => to_slv(opcode_type, 16#09#),
      1355 => to_slv(opcode_type, 16#11#),
      1356 => to_slv(opcode_type, 16#0B#),
      1357 => to_slv(opcode_type, 16#08#),
      1358 => to_slv(opcode_type, 16#0C#),
      1359 => to_slv(opcode_type, 16#30#),
      1360 => to_slv(opcode_type, 16#09#),
      1361 => to_slv(opcode_type, 16#08#),
      1362 => to_slv(opcode_type, 16#06#),
      1363 => to_slv(opcode_type, 16#0E#),
      1364 => to_slv(opcode_type, 16#9F#),
      1365 => to_slv(opcode_type, 16#08#),
      1366 => to_slv(opcode_type, 16#0B#),
      1367 => to_slv(opcode_type, 16#0A#),
      1368 => to_slv(opcode_type, 16#07#),
      1369 => to_slv(opcode_type, 16#07#),
      1370 => to_slv(opcode_type, 16#0C#),
      1371 => to_slv(opcode_type, 16#0E#),
      1372 => to_slv(opcode_type, 16#09#),
      1373 => to_slv(opcode_type, 16#0A#),
      1374 => to_slv(opcode_type, 16#95#),
      1375 to 1375 => (others => '0'),

      -- Program 43...
      1376 => to_slv(opcode_type, 16#09#),
      1377 => to_slv(opcode_type, 16#08#),
      1378 => to_slv(opcode_type, 16#08#),
      1379 => to_slv(opcode_type, 16#06#),
      1380 => to_slv(opcode_type, 16#11#),
      1381 => to_slv(opcode_type, 16#0C#),
      1382 => to_slv(opcode_type, 16#07#),
      1383 => to_slv(opcode_type, 16#0E#),
      1384 => to_slv(opcode_type, 16#0A#),
      1385 => to_slv(opcode_type, 16#08#),
      1386 => to_slv(opcode_type, 16#07#),
      1387 => to_slv(opcode_type, 16#0F#),
      1388 => to_slv(opcode_type, 16#0C#),
      1389 => to_slv(opcode_type, 16#08#),
      1390 => to_slv(opcode_type, 16#0E#),
      1391 => to_slv(opcode_type, 16#0E#),
      1392 => to_slv(opcode_type, 16#07#),
      1393 => to_slv(opcode_type, 16#08#),
      1394 => to_slv(opcode_type, 16#08#),
      1395 => to_slv(opcode_type, 16#0D#),
      1396 => to_slv(opcode_type, 16#26#),
      1397 => to_slv(opcode_type, 16#06#),
      1398 => to_slv(opcode_type, 16#0B#),
      1399 => to_slv(opcode_type, 16#98#),
      1400 => to_slv(opcode_type, 16#07#),
      1401 => to_slv(opcode_type, 16#07#),
      1402 => to_slv(opcode_type, 16#87#),
      1403 => to_slv(opcode_type, 16#0C#),
      1404 => to_slv(opcode_type, 16#09#),
      1405 => to_slv(opcode_type, 16#0A#),
      1406 => to_slv(opcode_type, 16#11#),
      1407 to 1407 => (others => '0'),

      -- Program 44...
      1408 => to_slv(opcode_type, 16#09#),
      1409 => to_slv(opcode_type, 16#07#),
      1410 => to_slv(opcode_type, 16#06#),
      1411 => to_slv(opcode_type, 16#06#),
      1412 => to_slv(opcode_type, 16#0D#),
      1413 => to_slv(opcode_type, 16#0C#),
      1414 => to_slv(opcode_type, 16#08#),
      1415 => to_slv(opcode_type, 16#A9#),
      1416 => to_slv(opcode_type, 16#0F#),
      1417 => to_slv(opcode_type, 16#06#),
      1418 => to_slv(opcode_type, 16#09#),
      1419 => to_slv(opcode_type, 16#0E#),
      1420 => to_slv(opcode_type, 16#0F#),
      1421 => to_slv(opcode_type, 16#09#),
      1422 => to_slv(opcode_type, 16#0A#),
      1423 => to_slv(opcode_type, 16#0F#),
      1424 => to_slv(opcode_type, 16#06#),
      1425 => to_slv(opcode_type, 16#08#),
      1426 => to_slv(opcode_type, 16#09#),
      1427 => to_slv(opcode_type, 16#0A#),
      1428 => to_slv(opcode_type, 16#0E#),
      1429 => to_slv(opcode_type, 16#09#),
      1430 => to_slv(opcode_type, 16#10#),
      1431 => to_slv(opcode_type, 16#0E#),
      1432 => to_slv(opcode_type, 16#09#),
      1433 => to_slv(opcode_type, 16#06#),
      1434 => to_slv(opcode_type, 16#9E#),
      1435 => to_slv(opcode_type, 16#10#),
      1436 => to_slv(opcode_type, 16#09#),
      1437 => to_slv(opcode_type, 16#0B#),
      1438 => to_slv(opcode_type, 16#FB#),
      1439 to 1439 => (others => '0'),

      -- Program 45...
      1440 => to_slv(opcode_type, 16#08#),
      1441 => to_slv(opcode_type, 16#06#),
      1442 => to_slv(opcode_type, 16#08#),
      1443 => to_slv(opcode_type, 16#08#),
      1444 => to_slv(opcode_type, 16#0B#),
      1445 => to_slv(opcode_type, 16#11#),
      1446 => to_slv(opcode_type, 16#06#),
      1447 => to_slv(opcode_type, 16#0B#),
      1448 => to_slv(opcode_type, 16#11#),
      1449 => to_slv(opcode_type, 16#06#),
      1450 => to_slv(opcode_type, 16#09#),
      1451 => to_slv(opcode_type, 16#0E#),
      1452 => to_slv(opcode_type, 16#0F#),
      1453 => to_slv(opcode_type, 16#08#),
      1454 => to_slv(opcode_type, 16#34#),
      1455 => to_slv(opcode_type, 16#38#),
      1456 => to_slv(opcode_type, 16#06#),
      1457 => to_slv(opcode_type, 16#06#),
      1458 => to_slv(opcode_type, 16#09#),
      1459 => to_slv(opcode_type, 16#11#),
      1460 => to_slv(opcode_type, 16#0B#),
      1461 => to_slv(opcode_type, 16#09#),
      1462 => to_slv(opcode_type, 16#0A#),
      1463 => to_slv(opcode_type, 16#0D#),
      1464 => to_slv(opcode_type, 16#09#),
      1465 => to_slv(opcode_type, 16#07#),
      1466 => to_slv(opcode_type, 16#0A#),
      1467 => to_slv(opcode_type, 16#0E#),
      1468 => to_slv(opcode_type, 16#08#),
      1469 => to_slv(opcode_type, 16#11#),
      1470 => to_slv(opcode_type, 16#0B#),
      1471 to 1471 => (others => '0'),

      -- Program 46...
      1472 => to_slv(opcode_type, 16#07#),
      1473 => to_slv(opcode_type, 16#09#),
      1474 => to_slv(opcode_type, 16#08#),
      1475 => to_slv(opcode_type, 16#08#),
      1476 => to_slv(opcode_type, 16#0D#),
      1477 => to_slv(opcode_type, 16#0D#),
      1478 => to_slv(opcode_type, 16#06#),
      1479 => to_slv(opcode_type, 16#0C#),
      1480 => to_slv(opcode_type, 16#0F#),
      1481 => to_slv(opcode_type, 16#07#),
      1482 => to_slv(opcode_type, 16#09#),
      1483 => to_slv(opcode_type, 16#0F#),
      1484 => to_slv(opcode_type, 16#11#),
      1485 => to_slv(opcode_type, 16#06#),
      1486 => to_slv(opcode_type, 16#0E#),
      1487 => to_slv(opcode_type, 16#11#),
      1488 => to_slv(opcode_type, 16#09#),
      1489 => to_slv(opcode_type, 16#07#),
      1490 => to_slv(opcode_type, 16#08#),
      1491 => to_slv(opcode_type, 16#0A#),
      1492 => to_slv(opcode_type, 16#0A#),
      1493 => to_slv(opcode_type, 16#09#),
      1494 => to_slv(opcode_type, 16#10#),
      1495 => to_slv(opcode_type, 16#0F#),
      1496 => to_slv(opcode_type, 16#08#),
      1497 => to_slv(opcode_type, 16#06#),
      1498 => to_slv(opcode_type, 16#0F#),
      1499 => to_slv(opcode_type, 16#10#),
      1500 => to_slv(opcode_type, 16#06#),
      1501 => to_slv(opcode_type, 16#10#),
      1502 => to_slv(opcode_type, 16#0F#),
      1503 to 1503 => (others => '0'),

      -- Program 47...
      1504 => to_slv(opcode_type, 16#09#),
      1505 => to_slv(opcode_type, 16#08#),
      1506 => to_slv(opcode_type, 16#09#),
      1507 => to_slv(opcode_type, 16#07#),
      1508 => to_slv(opcode_type, 16#0D#),
      1509 => to_slv(opcode_type, 16#0C#),
      1510 => to_slv(opcode_type, 16#09#),
      1511 => to_slv(opcode_type, 16#0B#),
      1512 => to_slv(opcode_type, 16#0E#),
      1513 => to_slv(opcode_type, 16#09#),
      1514 => to_slv(opcode_type, 16#07#),
      1515 => to_slv(opcode_type, 16#11#),
      1516 => to_slv(opcode_type, 16#91#),
      1517 => to_slv(opcode_type, 16#08#),
      1518 => to_slv(opcode_type, 16#0E#),
      1519 => to_slv(opcode_type, 16#0E#),
      1520 => to_slv(opcode_type, 16#09#),
      1521 => to_slv(opcode_type, 16#08#),
      1522 => to_slv(opcode_type, 16#08#),
      1523 => to_slv(opcode_type, 16#0A#),
      1524 => to_slv(opcode_type, 16#0B#),
      1525 => to_slv(opcode_type, 16#08#),
      1526 => to_slv(opcode_type, 16#A7#),
      1527 => to_slv(opcode_type, 16#0D#),
      1528 => to_slv(opcode_type, 16#08#),
      1529 => to_slv(opcode_type, 16#08#),
      1530 => to_slv(opcode_type, 16#0A#),
      1531 => to_slv(opcode_type, 16#0E#),
      1532 => to_slv(opcode_type, 16#09#),
      1533 => to_slv(opcode_type, 16#10#),
      1534 => to_slv(opcode_type, 16#0F#),
      1535 to 1535 => (others => '0'),

      -- Program 48...
      1536 => to_slv(opcode_type, 16#08#),
      1537 => to_slv(opcode_type, 16#09#),
      1538 => to_slv(opcode_type, 16#07#),
      1539 => to_slv(opcode_type, 16#07#),
      1540 => to_slv(opcode_type, 16#0D#),
      1541 => to_slv(opcode_type, 16#0B#),
      1542 => to_slv(opcode_type, 16#09#),
      1543 => to_slv(opcode_type, 16#11#),
      1544 => to_slv(opcode_type, 16#0A#),
      1545 => to_slv(opcode_type, 16#08#),
      1546 => to_slv(opcode_type, 16#08#),
      1547 => to_slv(opcode_type, 16#0B#),
      1548 => to_slv(opcode_type, 16#0E#),
      1549 => to_slv(opcode_type, 16#09#),
      1550 => to_slv(opcode_type, 16#BE#),
      1551 => to_slv(opcode_type, 16#0F#),
      1552 => to_slv(opcode_type, 16#08#),
      1553 => to_slv(opcode_type, 16#07#),
      1554 => to_slv(opcode_type, 16#07#),
      1555 => to_slv(opcode_type, 16#A5#),
      1556 => to_slv(opcode_type, 16#0D#),
      1557 => to_slv(opcode_type, 16#06#),
      1558 => to_slv(opcode_type, 16#10#),
      1559 => to_slv(opcode_type, 16#0F#),
      1560 => to_slv(opcode_type, 16#07#),
      1561 => to_slv(opcode_type, 16#06#),
      1562 => to_slv(opcode_type, 16#0C#),
      1563 => to_slv(opcode_type, 16#10#),
      1564 => to_slv(opcode_type, 16#07#),
      1565 => to_slv(opcode_type, 16#64#),
      1566 => to_slv(opcode_type, 16#0D#),
      1567 to 1567 => (others => '0'),

      -- Program 49...
      1568 => to_slv(opcode_type, 16#07#),
      1569 => to_slv(opcode_type, 16#09#),
      1570 => to_slv(opcode_type, 16#09#),
      1571 => to_slv(opcode_type, 16#07#),
      1572 => to_slv(opcode_type, 16#0F#),
      1573 => to_slv(opcode_type, 16#11#),
      1574 => to_slv(opcode_type, 16#08#),
      1575 => to_slv(opcode_type, 16#0B#),
      1576 => to_slv(opcode_type, 16#0D#),
      1577 => to_slv(opcode_type, 16#09#),
      1578 => to_slv(opcode_type, 16#06#),
      1579 => to_slv(opcode_type, 16#0D#),
      1580 => to_slv(opcode_type, 16#0A#),
      1581 => to_slv(opcode_type, 16#06#),
      1582 => to_slv(opcode_type, 16#CA#),
      1583 => to_slv(opcode_type, 16#0C#),
      1584 => to_slv(opcode_type, 16#06#),
      1585 => to_slv(opcode_type, 16#06#),
      1586 => to_slv(opcode_type, 16#09#),
      1587 => to_slv(opcode_type, 16#0B#),
      1588 => to_slv(opcode_type, 16#0D#),
      1589 => to_slv(opcode_type, 16#07#),
      1590 => to_slv(opcode_type, 16#0E#),
      1591 => to_slv(opcode_type, 16#0D#),
      1592 => to_slv(opcode_type, 16#06#),
      1593 => to_slv(opcode_type, 16#09#),
      1594 => to_slv(opcode_type, 16#EF#),
      1595 => to_slv(opcode_type, 16#0F#),
      1596 => to_slv(opcode_type, 16#09#),
      1597 => to_slv(opcode_type, 16#0F#),
      1598 => to_slv(opcode_type, 16#0C#),
      1599 to 1599 => (others => '0'),

      -- Program 50...
      1600 => to_slv(opcode_type, 16#06#),
      1601 => to_slv(opcode_type, 16#06#),
      1602 => to_slv(opcode_type, 16#06#),
      1603 => to_slv(opcode_type, 16#08#),
      1604 => to_slv(opcode_type, 16#0F#),
      1605 => to_slv(opcode_type, 16#0D#),
      1606 => to_slv(opcode_type, 16#06#),
      1607 => to_slv(opcode_type, 16#11#),
      1608 => to_slv(opcode_type, 16#11#),
      1609 => to_slv(opcode_type, 16#09#),
      1610 => to_slv(opcode_type, 16#08#),
      1611 => to_slv(opcode_type, 16#0D#),
      1612 => to_slv(opcode_type, 16#11#),
      1613 => to_slv(opcode_type, 16#07#),
      1614 => to_slv(opcode_type, 16#0E#),
      1615 => to_slv(opcode_type, 16#11#),
      1616 => to_slv(opcode_type, 16#08#),
      1617 => to_slv(opcode_type, 16#09#),
      1618 => to_slv(opcode_type, 16#08#),
      1619 => to_slv(opcode_type, 16#CE#),
      1620 => to_slv(opcode_type, 16#10#),
      1621 => to_slv(opcode_type, 16#06#),
      1622 => to_slv(opcode_type, 16#0D#),
      1623 => to_slv(opcode_type, 16#0A#),
      1624 => to_slv(opcode_type, 16#06#),
      1625 => to_slv(opcode_type, 16#07#),
      1626 => to_slv(opcode_type, 16#11#),
      1627 => to_slv(opcode_type, 16#30#),
      1628 => to_slv(opcode_type, 16#06#),
      1629 => to_slv(opcode_type, 16#0D#),
      1630 => to_slv(opcode_type, 16#D7#),
      1631 to 1631 => (others => '0'),

      -- Program 51...
      1632 => to_slv(opcode_type, 16#06#),
      1633 => to_slv(opcode_type, 16#07#),
      1634 => to_slv(opcode_type, 16#08#),
      1635 => to_slv(opcode_type, 16#06#),
      1636 => to_slv(opcode_type, 16#0E#),
      1637 => to_slv(opcode_type, 16#15#),
      1638 => to_slv(opcode_type, 16#06#),
      1639 => to_slv(opcode_type, 16#0A#),
      1640 => to_slv(opcode_type, 16#0F#),
      1641 => to_slv(opcode_type, 16#07#),
      1642 => to_slv(opcode_type, 16#08#),
      1643 => to_slv(opcode_type, 16#0E#),
      1644 => to_slv(opcode_type, 16#0B#),
      1645 => to_slv(opcode_type, 16#06#),
      1646 => to_slv(opcode_type, 16#10#),
      1647 => to_slv(opcode_type, 16#0B#),
      1648 => to_slv(opcode_type, 16#09#),
      1649 => to_slv(opcode_type, 16#08#),
      1650 => to_slv(opcode_type, 16#06#),
      1651 => to_slv(opcode_type, 16#10#),
      1652 => to_slv(opcode_type, 16#10#),
      1653 => to_slv(opcode_type, 16#09#),
      1654 => to_slv(opcode_type, 16#0A#),
      1655 => to_slv(opcode_type, 16#0C#),
      1656 => to_slv(opcode_type, 16#06#),
      1657 => to_slv(opcode_type, 16#09#),
      1658 => to_slv(opcode_type, 16#0E#),
      1659 => to_slv(opcode_type, 16#10#),
      1660 => to_slv(opcode_type, 16#06#),
      1661 => to_slv(opcode_type, 16#0D#),
      1662 => to_slv(opcode_type, 16#11#),
      1663 to 1663 => (others => '0'),

      -- Program 52...
      1664 => to_slv(opcode_type, 16#07#),
      1665 => to_slv(opcode_type, 16#06#),
      1666 => to_slv(opcode_type, 16#06#),
      1667 => to_slv(opcode_type, 16#09#),
      1668 => to_slv(opcode_type, 16#0B#),
      1669 => to_slv(opcode_type, 16#4B#),
      1670 => to_slv(opcode_type, 16#08#),
      1671 => to_slv(opcode_type, 16#10#),
      1672 => to_slv(opcode_type, 16#E0#),
      1673 => to_slv(opcode_type, 16#06#),
      1674 => to_slv(opcode_type, 16#08#),
      1675 => to_slv(opcode_type, 16#0A#),
      1676 => to_slv(opcode_type, 16#0A#),
      1677 => to_slv(opcode_type, 16#09#),
      1678 => to_slv(opcode_type, 16#11#),
      1679 => to_slv(opcode_type, 16#11#),
      1680 => to_slv(opcode_type, 16#07#),
      1681 => to_slv(opcode_type, 16#06#),
      1682 => to_slv(opcode_type, 16#07#),
      1683 => to_slv(opcode_type, 16#0B#),
      1684 => to_slv(opcode_type, 16#0B#),
      1685 => to_slv(opcode_type, 16#06#),
      1686 => to_slv(opcode_type, 16#0D#),
      1687 => to_slv(opcode_type, 16#0E#),
      1688 => to_slv(opcode_type, 16#08#),
      1689 => to_slv(opcode_type, 16#07#),
      1690 => to_slv(opcode_type, 16#11#),
      1691 => to_slv(opcode_type, 16#0D#),
      1692 => to_slv(opcode_type, 16#07#),
      1693 => to_slv(opcode_type, 16#0D#),
      1694 => to_slv(opcode_type, 16#10#),
      1695 to 1695 => (others => '0'),

      -- Program 53...
      1696 => to_slv(opcode_type, 16#07#),
      1697 => to_slv(opcode_type, 16#06#),
      1698 => to_slv(opcode_type, 16#09#),
      1699 => to_slv(opcode_type, 16#08#),
      1700 => to_slv(opcode_type, 16#0B#),
      1701 => to_slv(opcode_type, 16#11#),
      1702 => to_slv(opcode_type, 16#07#),
      1703 => to_slv(opcode_type, 16#0A#),
      1704 => to_slv(opcode_type, 16#0D#),
      1705 => to_slv(opcode_type, 16#09#),
      1706 => to_slv(opcode_type, 16#06#),
      1707 => to_slv(opcode_type, 16#0B#),
      1708 => to_slv(opcode_type, 16#10#),
      1709 => to_slv(opcode_type, 16#06#),
      1710 => to_slv(opcode_type, 16#11#),
      1711 => to_slv(opcode_type, 16#FF#),
      1712 => to_slv(opcode_type, 16#09#),
      1713 => to_slv(opcode_type, 16#08#),
      1714 => to_slv(opcode_type, 16#08#),
      1715 => to_slv(opcode_type, 16#0F#),
      1716 => to_slv(opcode_type, 16#0D#),
      1717 => to_slv(opcode_type, 16#09#),
      1718 => to_slv(opcode_type, 16#0B#),
      1719 => to_slv(opcode_type, 16#0C#),
      1720 => to_slv(opcode_type, 16#06#),
      1721 => to_slv(opcode_type, 16#08#),
      1722 => to_slv(opcode_type, 16#0B#),
      1723 => to_slv(opcode_type, 16#0F#),
      1724 => to_slv(opcode_type, 16#06#),
      1725 => to_slv(opcode_type, 16#11#),
      1726 => to_slv(opcode_type, 16#0C#),
      1727 to 1727 => (others => '0'),

      -- Program 54...
      1728 => to_slv(opcode_type, 16#08#),
      1729 => to_slv(opcode_type, 16#06#),
      1730 => to_slv(opcode_type, 16#08#),
      1731 => to_slv(opcode_type, 16#08#),
      1732 => to_slv(opcode_type, 16#10#),
      1733 => to_slv(opcode_type, 16#0D#),
      1734 => to_slv(opcode_type, 16#08#),
      1735 => to_slv(opcode_type, 16#0F#),
      1736 => to_slv(opcode_type, 16#8D#),
      1737 => to_slv(opcode_type, 16#08#),
      1738 => to_slv(opcode_type, 16#06#),
      1739 => to_slv(opcode_type, 16#0F#),
      1740 => to_slv(opcode_type, 16#10#),
      1741 => to_slv(opcode_type, 16#09#),
      1742 => to_slv(opcode_type, 16#11#),
      1743 => to_slv(opcode_type, 16#0B#),
      1744 => to_slv(opcode_type, 16#07#),
      1745 => to_slv(opcode_type, 16#08#),
      1746 => to_slv(opcode_type, 16#08#),
      1747 => to_slv(opcode_type, 16#0D#),
      1748 => to_slv(opcode_type, 16#10#),
      1749 => to_slv(opcode_type, 16#06#),
      1750 => to_slv(opcode_type, 16#10#),
      1751 => to_slv(opcode_type, 16#0D#),
      1752 => to_slv(opcode_type, 16#08#),
      1753 => to_slv(opcode_type, 16#07#),
      1754 => to_slv(opcode_type, 16#0C#),
      1755 => to_slv(opcode_type, 16#0E#),
      1756 => to_slv(opcode_type, 16#07#),
      1757 => to_slv(opcode_type, 16#0E#),
      1758 => to_slv(opcode_type, 16#0F#),
      1759 to 1759 => (others => '0'),

      -- Program 55...
      1760 => to_slv(opcode_type, 16#09#),
      1761 => to_slv(opcode_type, 16#09#),
      1762 => to_slv(opcode_type, 16#09#),
      1763 => to_slv(opcode_type, 16#08#),
      1764 => to_slv(opcode_type, 16#0B#),
      1765 => to_slv(opcode_type, 16#10#),
      1766 => to_slv(opcode_type, 16#06#),
      1767 => to_slv(opcode_type, 16#0E#),
      1768 => to_slv(opcode_type, 16#11#),
      1769 => to_slv(opcode_type, 16#07#),
      1770 => to_slv(opcode_type, 16#08#),
      1771 => to_slv(opcode_type, 16#10#),
      1772 => to_slv(opcode_type, 16#10#),
      1773 => to_slv(opcode_type, 16#07#),
      1774 => to_slv(opcode_type, 16#0C#),
      1775 => to_slv(opcode_type, 16#11#),
      1776 => to_slv(opcode_type, 16#07#),
      1777 => to_slv(opcode_type, 16#06#),
      1778 => to_slv(opcode_type, 16#07#),
      1779 => to_slv(opcode_type, 16#0C#),
      1780 => to_slv(opcode_type, 16#0F#),
      1781 => to_slv(opcode_type, 16#07#),
      1782 => to_slv(opcode_type, 16#E2#),
      1783 => to_slv(opcode_type, 16#0A#),
      1784 => to_slv(opcode_type, 16#07#),
      1785 => to_slv(opcode_type, 16#07#),
      1786 => to_slv(opcode_type, 16#0B#),
      1787 => to_slv(opcode_type, 16#0B#),
      1788 => to_slv(opcode_type, 16#08#),
      1789 => to_slv(opcode_type, 16#33#),
      1790 => to_slv(opcode_type, 16#0D#),
      1791 to 1791 => (others => '0'),

      -- Program 56...
      1792 => to_slv(opcode_type, 16#07#),
      1793 => to_slv(opcode_type, 16#06#),
      1794 => to_slv(opcode_type, 16#07#),
      1795 => to_slv(opcode_type, 16#09#),
      1796 => to_slv(opcode_type, 16#10#),
      1797 => to_slv(opcode_type, 16#10#),
      1798 => to_slv(opcode_type, 16#07#),
      1799 => to_slv(opcode_type, 16#0C#),
      1800 => to_slv(opcode_type, 16#0E#),
      1801 => to_slv(opcode_type, 16#06#),
      1802 => to_slv(opcode_type, 16#09#),
      1803 => to_slv(opcode_type, 16#0D#),
      1804 => to_slv(opcode_type, 16#0A#),
      1805 => to_slv(opcode_type, 16#09#),
      1806 => to_slv(opcode_type, 16#0A#),
      1807 => to_slv(opcode_type, 16#0F#),
      1808 => to_slv(opcode_type, 16#09#),
      1809 => to_slv(opcode_type, 16#08#),
      1810 => to_slv(opcode_type, 16#06#),
      1811 => to_slv(opcode_type, 16#10#),
      1812 => to_slv(opcode_type, 16#0C#),
      1813 => to_slv(opcode_type, 16#06#),
      1814 => to_slv(opcode_type, 16#0C#),
      1815 => to_slv(opcode_type, 16#11#),
      1816 => to_slv(opcode_type, 16#06#),
      1817 => to_slv(opcode_type, 16#08#),
      1818 => to_slv(opcode_type, 16#0F#),
      1819 => to_slv(opcode_type, 16#10#),
      1820 => to_slv(opcode_type, 16#06#),
      1821 => to_slv(opcode_type, 16#95#),
      1822 => to_slv(opcode_type, 16#0F#),
      1823 to 1823 => (others => '0'),

      -- Program 57...
      1824 => to_slv(opcode_type, 16#09#),
      1825 => to_slv(opcode_type, 16#08#),
      1826 => to_slv(opcode_type, 16#07#),
      1827 => to_slv(opcode_type, 16#08#),
      1828 => to_slv(opcode_type, 16#10#),
      1829 => to_slv(opcode_type, 16#10#),
      1830 => to_slv(opcode_type, 16#08#),
      1831 => to_slv(opcode_type, 16#0E#),
      1832 => to_slv(opcode_type, 16#0A#),
      1833 => to_slv(opcode_type, 16#08#),
      1834 => to_slv(opcode_type, 16#07#),
      1835 => to_slv(opcode_type, 16#10#),
      1836 => to_slv(opcode_type, 16#0E#),
      1837 => to_slv(opcode_type, 16#08#),
      1838 => to_slv(opcode_type, 16#0D#),
      1839 => to_slv(opcode_type, 16#0F#),
      1840 => to_slv(opcode_type, 16#07#),
      1841 => to_slv(opcode_type, 16#09#),
      1842 => to_slv(opcode_type, 16#07#),
      1843 => to_slv(opcode_type, 16#11#),
      1844 => to_slv(opcode_type, 16#0D#),
      1845 => to_slv(opcode_type, 16#07#),
      1846 => to_slv(opcode_type, 16#0E#),
      1847 => to_slv(opcode_type, 16#0B#),
      1848 => to_slv(opcode_type, 16#08#),
      1849 => to_slv(opcode_type, 16#09#),
      1850 => to_slv(opcode_type, 16#0E#),
      1851 => to_slv(opcode_type, 16#2A#),
      1852 => to_slv(opcode_type, 16#07#),
      1853 => to_slv(opcode_type, 16#0E#),
      1854 => to_slv(opcode_type, 16#0F#),
      1855 to 1855 => (others => '0'),

      -- Program 58...
      1856 => to_slv(opcode_type, 16#09#),
      1857 => to_slv(opcode_type, 16#07#),
      1858 => to_slv(opcode_type, 16#07#),
      1859 => to_slv(opcode_type, 16#07#),
      1860 => to_slv(opcode_type, 16#0A#),
      1861 => to_slv(opcode_type, 16#0A#),
      1862 => to_slv(opcode_type, 16#07#),
      1863 => to_slv(opcode_type, 16#0E#),
      1864 => to_slv(opcode_type, 16#11#),
      1865 => to_slv(opcode_type, 16#08#),
      1866 => to_slv(opcode_type, 16#08#),
      1867 => to_slv(opcode_type, 16#D8#),
      1868 => to_slv(opcode_type, 16#0F#),
      1869 => to_slv(opcode_type, 16#08#),
      1870 => to_slv(opcode_type, 16#10#),
      1871 => to_slv(opcode_type, 16#0D#),
      1872 => to_slv(opcode_type, 16#08#),
      1873 => to_slv(opcode_type, 16#08#),
      1874 => to_slv(opcode_type, 16#07#),
      1875 => to_slv(opcode_type, 16#4F#),
      1876 => to_slv(opcode_type, 16#10#),
      1877 => to_slv(opcode_type, 16#06#),
      1878 => to_slv(opcode_type, 16#22#),
      1879 => to_slv(opcode_type, 16#11#),
      1880 => to_slv(opcode_type, 16#07#),
      1881 => to_slv(opcode_type, 16#07#),
      1882 => to_slv(opcode_type, 16#0C#),
      1883 => to_slv(opcode_type, 16#11#),
      1884 => to_slv(opcode_type, 16#08#),
      1885 => to_slv(opcode_type, 16#11#),
      1886 => to_slv(opcode_type, 16#0F#),
      1887 to 1887 => (others => '0'),

      -- Program 59...
      1888 => to_slv(opcode_type, 16#06#),
      1889 => to_slv(opcode_type, 16#06#),
      1890 => to_slv(opcode_type, 16#06#),
      1891 => to_slv(opcode_type, 16#07#),
      1892 => to_slv(opcode_type, 16#0D#),
      1893 => to_slv(opcode_type, 16#0A#),
      1894 => to_slv(opcode_type, 16#09#),
      1895 => to_slv(opcode_type, 16#0E#),
      1896 => to_slv(opcode_type, 16#0B#),
      1897 => to_slv(opcode_type, 16#09#),
      1898 => to_slv(opcode_type, 16#07#),
      1899 => to_slv(opcode_type, 16#0D#),
      1900 => to_slv(opcode_type, 16#0C#),
      1901 => to_slv(opcode_type, 16#06#),
      1902 => to_slv(opcode_type, 16#11#),
      1903 => to_slv(opcode_type, 16#10#),
      1904 => to_slv(opcode_type, 16#07#),
      1905 => to_slv(opcode_type, 16#08#),
      1906 => to_slv(opcode_type, 16#07#),
      1907 => to_slv(opcode_type, 16#0E#),
      1908 => to_slv(opcode_type, 16#0A#),
      1909 => to_slv(opcode_type, 16#09#),
      1910 => to_slv(opcode_type, 16#0F#),
      1911 => to_slv(opcode_type, 16#11#),
      1912 => to_slv(opcode_type, 16#06#),
      1913 => to_slv(opcode_type, 16#09#),
      1914 => to_slv(opcode_type, 16#0A#),
      1915 => to_slv(opcode_type, 16#0B#),
      1916 => to_slv(opcode_type, 16#09#),
      1917 => to_slv(opcode_type, 16#0B#),
      1918 => to_slv(opcode_type, 16#B9#),
      1919 to 1919 => (others => '0'),

      -- Program 60...
      1920 => to_slv(opcode_type, 16#08#),
      1921 => to_slv(opcode_type, 16#07#),
      1922 => to_slv(opcode_type, 16#06#),
      1923 => to_slv(opcode_type, 16#07#),
      1924 => to_slv(opcode_type, 16#0E#),
      1925 => to_slv(opcode_type, 16#0B#),
      1926 => to_slv(opcode_type, 16#06#),
      1927 => to_slv(opcode_type, 16#10#),
      1928 => to_slv(opcode_type, 16#0B#),
      1929 => to_slv(opcode_type, 16#07#),
      1930 => to_slv(opcode_type, 16#09#),
      1931 => to_slv(opcode_type, 16#0D#),
      1932 => to_slv(opcode_type, 16#0C#),
      1933 => to_slv(opcode_type, 16#08#),
      1934 => to_slv(opcode_type, 16#0F#),
      1935 => to_slv(opcode_type, 16#11#),
      1936 => to_slv(opcode_type, 16#06#),
      1937 => to_slv(opcode_type, 16#07#),
      1938 => to_slv(opcode_type, 16#09#),
      1939 => to_slv(opcode_type, 16#51#),
      1940 => to_slv(opcode_type, 16#0E#),
      1941 => to_slv(opcode_type, 16#07#),
      1942 => to_slv(opcode_type, 16#0D#),
      1943 => to_slv(opcode_type, 16#0C#),
      1944 => to_slv(opcode_type, 16#06#),
      1945 => to_slv(opcode_type, 16#07#),
      1946 => to_slv(opcode_type, 16#10#),
      1947 => to_slv(opcode_type, 16#0A#),
      1948 => to_slv(opcode_type, 16#07#),
      1949 => to_slv(opcode_type, 16#0B#),
      1950 => to_slv(opcode_type, 16#91#),
      1951 to 1951 => (others => '0'),

      -- Program 61...
      1952 => to_slv(opcode_type, 16#06#),
      1953 => to_slv(opcode_type, 16#06#),
      1954 => to_slv(opcode_type, 16#07#),
      1955 => to_slv(opcode_type, 16#07#),
      1956 => to_slv(opcode_type, 16#11#),
      1957 => to_slv(opcode_type, 16#10#),
      1958 => to_slv(opcode_type, 16#09#),
      1959 => to_slv(opcode_type, 16#0A#),
      1960 => to_slv(opcode_type, 16#0D#),
      1961 => to_slv(opcode_type, 16#06#),
      1962 => to_slv(opcode_type, 16#07#),
      1963 => to_slv(opcode_type, 16#10#),
      1964 => to_slv(opcode_type, 16#0E#),
      1965 => to_slv(opcode_type, 16#09#),
      1966 => to_slv(opcode_type, 16#11#),
      1967 => to_slv(opcode_type, 16#0C#),
      1968 => to_slv(opcode_type, 16#06#),
      1969 => to_slv(opcode_type, 16#07#),
      1970 => to_slv(opcode_type, 16#07#),
      1971 => to_slv(opcode_type, 16#10#),
      1972 => to_slv(opcode_type, 16#0C#),
      1973 => to_slv(opcode_type, 16#06#),
      1974 => to_slv(opcode_type, 16#0F#),
      1975 => to_slv(opcode_type, 16#0E#),
      1976 => to_slv(opcode_type, 16#06#),
      1977 => to_slv(opcode_type, 16#08#),
      1978 => to_slv(opcode_type, 16#10#),
      1979 => to_slv(opcode_type, 16#10#),
      1980 => to_slv(opcode_type, 16#09#),
      1981 => to_slv(opcode_type, 16#0B#),
      1982 => to_slv(opcode_type, 16#0C#),
      1983 to 1983 => (others => '0'),

      -- Program 62...
      1984 => to_slv(opcode_type, 16#08#),
      1985 => to_slv(opcode_type, 16#08#),
      1986 => to_slv(opcode_type, 16#06#),
      1987 => to_slv(opcode_type, 16#07#),
      1988 => to_slv(opcode_type, 16#98#),
      1989 => to_slv(opcode_type, 16#0C#),
      1990 => to_slv(opcode_type, 16#09#),
      1991 => to_slv(opcode_type, 16#0B#),
      1992 => to_slv(opcode_type, 16#0A#),
      1993 => to_slv(opcode_type, 16#08#),
      1994 => to_slv(opcode_type, 16#09#),
      1995 => to_slv(opcode_type, 16#36#),
      1996 => to_slv(opcode_type, 16#11#),
      1997 => to_slv(opcode_type, 16#09#),
      1998 => to_slv(opcode_type, 16#0E#),
      1999 => to_slv(opcode_type, 16#0E#),
      2000 => to_slv(opcode_type, 16#06#),
      2001 => to_slv(opcode_type, 16#09#),
      2002 => to_slv(opcode_type, 16#08#),
      2003 => to_slv(opcode_type, 16#0D#),
      2004 => to_slv(opcode_type, 16#0C#),
      2005 => to_slv(opcode_type, 16#07#),
      2006 => to_slv(opcode_type, 16#0D#),
      2007 => to_slv(opcode_type, 16#11#),
      2008 => to_slv(opcode_type, 16#06#),
      2009 => to_slv(opcode_type, 16#07#),
      2010 => to_slv(opcode_type, 16#0E#),
      2011 => to_slv(opcode_type, 16#D3#),
      2012 => to_slv(opcode_type, 16#08#),
      2013 => to_slv(opcode_type, 16#0E#),
      2014 => to_slv(opcode_type, 16#F9#),
      2015 to 2015 => (others => '0'),

      -- Program 63...
      2016 => to_slv(opcode_type, 16#08#),
      2017 => to_slv(opcode_type, 16#09#),
      2018 => to_slv(opcode_type, 16#08#),
      2019 => to_slv(opcode_type, 16#07#),
      2020 => to_slv(opcode_type, 16#0D#),
      2021 => to_slv(opcode_type, 16#0C#),
      2022 => to_slv(opcode_type, 16#07#),
      2023 => to_slv(opcode_type, 16#0F#),
      2024 => to_slv(opcode_type, 16#0F#),
      2025 => to_slv(opcode_type, 16#06#),
      2026 => to_slv(opcode_type, 16#09#),
      2027 => to_slv(opcode_type, 16#0C#),
      2028 => to_slv(opcode_type, 16#0F#),
      2029 => to_slv(opcode_type, 16#07#),
      2030 => to_slv(opcode_type, 16#0E#),
      2031 => to_slv(opcode_type, 16#11#),
      2032 => to_slv(opcode_type, 16#07#),
      2033 => to_slv(opcode_type, 16#06#),
      2034 => to_slv(opcode_type, 16#08#),
      2035 => to_slv(opcode_type, 16#0B#),
      2036 => to_slv(opcode_type, 16#10#),
      2037 => to_slv(opcode_type, 16#09#),
      2038 => to_slv(opcode_type, 16#0B#),
      2039 => to_slv(opcode_type, 16#10#),
      2040 => to_slv(opcode_type, 16#08#),
      2041 => to_slv(opcode_type, 16#08#),
      2042 => to_slv(opcode_type, 16#11#),
      2043 => to_slv(opcode_type, 16#0F#),
      2044 => to_slv(opcode_type, 16#07#),
      2045 => to_slv(opcode_type, 16#0A#),
      2046 => to_slv(opcode_type, 16#0A#),
      2047 to 2047 => (others => '0'),

      -- Program 64...
      2048 => to_slv(opcode_type, 16#06#),
      2049 => to_slv(opcode_type, 16#07#),
      2050 => to_slv(opcode_type, 16#09#),
      2051 => to_slv(opcode_type, 16#08#),
      2052 => to_slv(opcode_type, 16#11#),
      2053 => to_slv(opcode_type, 16#0F#),
      2054 => to_slv(opcode_type, 16#07#),
      2055 => to_slv(opcode_type, 16#0B#),
      2056 => to_slv(opcode_type, 16#0F#),
      2057 => to_slv(opcode_type, 16#07#),
      2058 => to_slv(opcode_type, 16#08#),
      2059 => to_slv(opcode_type, 16#11#),
      2060 => to_slv(opcode_type, 16#0D#),
      2061 => to_slv(opcode_type, 16#06#),
      2062 => to_slv(opcode_type, 16#0C#),
      2063 => to_slv(opcode_type, 16#0F#),
      2064 => to_slv(opcode_type, 16#09#),
      2065 => to_slv(opcode_type, 16#08#),
      2066 => to_slv(opcode_type, 16#07#),
      2067 => to_slv(opcode_type, 16#10#),
      2068 => to_slv(opcode_type, 16#0A#),
      2069 => to_slv(opcode_type, 16#08#),
      2070 => to_slv(opcode_type, 16#0A#),
      2071 => to_slv(opcode_type, 16#0F#),
      2072 => to_slv(opcode_type, 16#08#),
      2073 => to_slv(opcode_type, 16#07#),
      2074 => to_slv(opcode_type, 16#0F#),
      2075 => to_slv(opcode_type, 16#0E#),
      2076 => to_slv(opcode_type, 16#09#),
      2077 => to_slv(opcode_type, 16#0D#),
      2078 => to_slv(opcode_type, 16#0F#),
      2079 to 2079 => (others => '0'),

      -- Program 65...
      2080 => to_slv(opcode_type, 16#07#),
      2081 => to_slv(opcode_type, 16#09#),
      2082 => to_slv(opcode_type, 16#08#),
      2083 => to_slv(opcode_type, 16#07#),
      2084 => to_slv(opcode_type, 16#0F#),
      2085 => to_slv(opcode_type, 16#0E#),
      2086 => to_slv(opcode_type, 16#09#),
      2087 => to_slv(opcode_type, 16#0E#),
      2088 => to_slv(opcode_type, 16#10#),
      2089 => to_slv(opcode_type, 16#08#),
      2090 => to_slv(opcode_type, 16#07#),
      2091 => to_slv(opcode_type, 16#0E#),
      2092 => to_slv(opcode_type, 16#0F#),
      2093 => to_slv(opcode_type, 16#07#),
      2094 => to_slv(opcode_type, 16#0B#),
      2095 => to_slv(opcode_type, 16#10#),
      2096 => to_slv(opcode_type, 16#08#),
      2097 => to_slv(opcode_type, 16#07#),
      2098 => to_slv(opcode_type, 16#07#),
      2099 => to_slv(opcode_type, 16#11#),
      2100 => to_slv(opcode_type, 16#0E#),
      2101 => to_slv(opcode_type, 16#07#),
      2102 => to_slv(opcode_type, 16#10#),
      2103 => to_slv(opcode_type, 16#0D#),
      2104 => to_slv(opcode_type, 16#07#),
      2105 => to_slv(opcode_type, 16#09#),
      2106 => to_slv(opcode_type, 16#0E#),
      2107 => to_slv(opcode_type, 16#0E#),
      2108 => to_slv(opcode_type, 16#07#),
      2109 => to_slv(opcode_type, 16#0D#),
      2110 => to_slv(opcode_type, 16#0C#),
      2111 to 2111 => (others => '0'),

      -- Program 66...
      2112 => to_slv(opcode_type, 16#08#),
      2113 => to_slv(opcode_type, 16#07#),
      2114 => to_slv(opcode_type, 16#09#),
      2115 => to_slv(opcode_type, 16#08#),
      2116 => to_slv(opcode_type, 16#0E#),
      2117 => to_slv(opcode_type, 16#0A#),
      2118 => to_slv(opcode_type, 16#08#),
      2119 => to_slv(opcode_type, 16#0C#),
      2120 => to_slv(opcode_type, 16#10#),
      2121 => to_slv(opcode_type, 16#08#),
      2122 => to_slv(opcode_type, 16#09#),
      2123 => to_slv(opcode_type, 16#0F#),
      2124 => to_slv(opcode_type, 16#0E#),
      2125 => to_slv(opcode_type, 16#06#),
      2126 => to_slv(opcode_type, 16#9B#),
      2127 => to_slv(opcode_type, 16#0C#),
      2128 => to_slv(opcode_type, 16#06#),
      2129 => to_slv(opcode_type, 16#08#),
      2130 => to_slv(opcode_type, 16#08#),
      2131 => to_slv(opcode_type, 16#0A#),
      2132 => to_slv(opcode_type, 16#0E#),
      2133 => to_slv(opcode_type, 16#06#),
      2134 => to_slv(opcode_type, 16#0B#),
      2135 => to_slv(opcode_type, 16#0D#),
      2136 => to_slv(opcode_type, 16#07#),
      2137 => to_slv(opcode_type, 16#07#),
      2138 => to_slv(opcode_type, 16#0A#),
      2139 => to_slv(opcode_type, 16#0E#),
      2140 => to_slv(opcode_type, 16#09#),
      2141 => to_slv(opcode_type, 16#9F#),
      2142 => to_slv(opcode_type, 16#10#),
      2143 to 2143 => (others => '0'),

      -- Program 67...
      2144 => to_slv(opcode_type, 16#09#),
      2145 => to_slv(opcode_type, 16#09#),
      2146 => to_slv(opcode_type, 16#08#),
      2147 => to_slv(opcode_type, 16#09#),
      2148 => to_slv(opcode_type, 16#0C#),
      2149 => to_slv(opcode_type, 16#0B#),
      2150 => to_slv(opcode_type, 16#07#),
      2151 => to_slv(opcode_type, 16#54#),
      2152 => to_slv(opcode_type, 16#0F#),
      2153 => to_slv(opcode_type, 16#06#),
      2154 => to_slv(opcode_type, 16#09#),
      2155 => to_slv(opcode_type, 16#0D#),
      2156 => to_slv(opcode_type, 16#0A#),
      2157 => to_slv(opcode_type, 16#09#),
      2158 => to_slv(opcode_type, 16#0B#),
      2159 => to_slv(opcode_type, 16#0E#),
      2160 => to_slv(opcode_type, 16#07#),
      2161 => to_slv(opcode_type, 16#08#),
      2162 => to_slv(opcode_type, 16#06#),
      2163 => to_slv(opcode_type, 16#10#),
      2164 => to_slv(opcode_type, 16#0E#),
      2165 => to_slv(opcode_type, 16#09#),
      2166 => to_slv(opcode_type, 16#0C#),
      2167 => to_slv(opcode_type, 16#11#),
      2168 => to_slv(opcode_type, 16#08#),
      2169 => to_slv(opcode_type, 16#09#),
      2170 => to_slv(opcode_type, 16#0E#),
      2171 => to_slv(opcode_type, 16#0A#),
      2172 => to_slv(opcode_type, 16#08#),
      2173 => to_slv(opcode_type, 16#0E#),
      2174 => to_slv(opcode_type, 16#10#),
      2175 to 2175 => (others => '0'),

      -- Program 68...
      2176 => to_slv(opcode_type, 16#08#),
      2177 => to_slv(opcode_type, 16#09#),
      2178 => to_slv(opcode_type, 16#09#),
      2179 => to_slv(opcode_type, 16#09#),
      2180 => to_slv(opcode_type, 16#0C#),
      2181 => to_slv(opcode_type, 16#0C#),
      2182 => to_slv(opcode_type, 16#06#),
      2183 => to_slv(opcode_type, 16#0F#),
      2184 => to_slv(opcode_type, 16#6C#),
      2185 => to_slv(opcode_type, 16#06#),
      2186 => to_slv(opcode_type, 16#09#),
      2187 => to_slv(opcode_type, 16#0A#),
      2188 => to_slv(opcode_type, 16#10#),
      2189 => to_slv(opcode_type, 16#09#),
      2190 => to_slv(opcode_type, 16#11#),
      2191 => to_slv(opcode_type, 16#0C#),
      2192 => to_slv(opcode_type, 16#06#),
      2193 => to_slv(opcode_type, 16#08#),
      2194 => to_slv(opcode_type, 16#08#),
      2195 => to_slv(opcode_type, 16#0E#),
      2196 => to_slv(opcode_type, 16#0A#),
      2197 => to_slv(opcode_type, 16#07#),
      2198 => to_slv(opcode_type, 16#11#),
      2199 => to_slv(opcode_type, 16#0E#),
      2200 => to_slv(opcode_type, 16#09#),
      2201 => to_slv(opcode_type, 16#06#),
      2202 => to_slv(opcode_type, 16#0D#),
      2203 => to_slv(opcode_type, 16#0D#),
      2204 => to_slv(opcode_type, 16#08#),
      2205 => to_slv(opcode_type, 16#10#),
      2206 => to_slv(opcode_type, 16#10#),
      2207 to 2207 => (others => '0'),

      -- Program 69...
      2208 => to_slv(opcode_type, 16#09#),
      2209 => to_slv(opcode_type, 16#09#),
      2210 => to_slv(opcode_type, 16#08#),
      2211 => to_slv(opcode_type, 16#07#),
      2212 => to_slv(opcode_type, 16#0A#),
      2213 => to_slv(opcode_type, 16#0F#),
      2214 => to_slv(opcode_type, 16#09#),
      2215 => to_slv(opcode_type, 16#0D#),
      2216 => to_slv(opcode_type, 16#71#),
      2217 => to_slv(opcode_type, 16#08#),
      2218 => to_slv(opcode_type, 16#06#),
      2219 => to_slv(opcode_type, 16#10#),
      2220 => to_slv(opcode_type, 16#0C#),
      2221 => to_slv(opcode_type, 16#07#),
      2222 => to_slv(opcode_type, 16#0F#),
      2223 => to_slv(opcode_type, 16#11#),
      2224 => to_slv(opcode_type, 16#08#),
      2225 => to_slv(opcode_type, 16#06#),
      2226 => to_slv(opcode_type, 16#06#),
      2227 => to_slv(opcode_type, 16#11#),
      2228 => to_slv(opcode_type, 16#0A#),
      2229 => to_slv(opcode_type, 16#06#),
      2230 => to_slv(opcode_type, 16#0B#),
      2231 => to_slv(opcode_type, 16#11#),
      2232 => to_slv(opcode_type, 16#06#),
      2233 => to_slv(opcode_type, 16#09#),
      2234 => to_slv(opcode_type, 16#0E#),
      2235 => to_slv(opcode_type, 16#0B#),
      2236 => to_slv(opcode_type, 16#06#),
      2237 => to_slv(opcode_type, 16#0D#),
      2238 => to_slv(opcode_type, 16#0A#),
      2239 to 2239 => (others => '0'),

      -- Program 70...
      2240 => to_slv(opcode_type, 16#06#),
      2241 => to_slv(opcode_type, 16#06#),
      2242 => to_slv(opcode_type, 16#06#),
      2243 => to_slv(opcode_type, 16#06#),
      2244 => to_slv(opcode_type, 16#4D#),
      2245 => to_slv(opcode_type, 16#11#),
      2246 => to_slv(opcode_type, 16#09#),
      2247 => to_slv(opcode_type, 16#0A#),
      2248 => to_slv(opcode_type, 16#0C#),
      2249 => to_slv(opcode_type, 16#09#),
      2250 => to_slv(opcode_type, 16#06#),
      2251 => to_slv(opcode_type, 16#0B#),
      2252 => to_slv(opcode_type, 16#0E#),
      2253 => to_slv(opcode_type, 16#09#),
      2254 => to_slv(opcode_type, 16#0B#),
      2255 => to_slv(opcode_type, 16#0D#),
      2256 => to_slv(opcode_type, 16#06#),
      2257 => to_slv(opcode_type, 16#06#),
      2258 => to_slv(opcode_type, 16#06#),
      2259 => to_slv(opcode_type, 16#0B#),
      2260 => to_slv(opcode_type, 16#11#),
      2261 => to_slv(opcode_type, 16#06#),
      2262 => to_slv(opcode_type, 16#10#),
      2263 => to_slv(opcode_type, 16#0F#),
      2264 => to_slv(opcode_type, 16#06#),
      2265 => to_slv(opcode_type, 16#09#),
      2266 => to_slv(opcode_type, 16#0F#),
      2267 => to_slv(opcode_type, 16#0B#),
      2268 => to_slv(opcode_type, 16#07#),
      2269 => to_slv(opcode_type, 16#0B#),
      2270 => to_slv(opcode_type, 16#0B#),
      2271 to 2271 => (others => '0'),

      -- Program 71...
      2272 => to_slv(opcode_type, 16#08#),
      2273 => to_slv(opcode_type, 16#09#),
      2274 => to_slv(opcode_type, 16#09#),
      2275 => to_slv(opcode_type, 16#08#),
      2276 => to_slv(opcode_type, 16#0A#),
      2277 => to_slv(opcode_type, 16#0F#),
      2278 => to_slv(opcode_type, 16#06#),
      2279 => to_slv(opcode_type, 16#10#),
      2280 => to_slv(opcode_type, 16#76#),
      2281 => to_slv(opcode_type, 16#09#),
      2282 => to_slv(opcode_type, 16#06#),
      2283 => to_slv(opcode_type, 16#0A#),
      2284 => to_slv(opcode_type, 16#10#),
      2285 => to_slv(opcode_type, 16#09#),
      2286 => to_slv(opcode_type, 16#10#),
      2287 => to_slv(opcode_type, 16#0E#),
      2288 => to_slv(opcode_type, 16#09#),
      2289 => to_slv(opcode_type, 16#07#),
      2290 => to_slv(opcode_type, 16#06#),
      2291 => to_slv(opcode_type, 16#0E#),
      2292 => to_slv(opcode_type, 16#10#),
      2293 => to_slv(opcode_type, 16#09#),
      2294 => to_slv(opcode_type, 16#11#),
      2295 => to_slv(opcode_type, 16#11#),
      2296 => to_slv(opcode_type, 16#09#),
      2297 => to_slv(opcode_type, 16#07#),
      2298 => to_slv(opcode_type, 16#0B#),
      2299 => to_slv(opcode_type, 16#0A#),
      2300 => to_slv(opcode_type, 16#09#),
      2301 => to_slv(opcode_type, 16#3E#),
      2302 => to_slv(opcode_type, 16#10#),
      2303 to 2303 => (others => '0'),

      -- Program 72...
      2304 => to_slv(opcode_type, 16#09#),
      2305 => to_slv(opcode_type, 16#08#),
      2306 => to_slv(opcode_type, 16#07#),
      2307 => to_slv(opcode_type, 16#09#),
      2308 => to_slv(opcode_type, 16#B6#),
      2309 => to_slv(opcode_type, 16#0B#),
      2310 => to_slv(opcode_type, 16#08#),
      2311 => to_slv(opcode_type, 16#0A#),
      2312 => to_slv(opcode_type, 16#0E#),
      2313 => to_slv(opcode_type, 16#09#),
      2314 => to_slv(opcode_type, 16#06#),
      2315 => to_slv(opcode_type, 16#10#),
      2316 => to_slv(opcode_type, 16#10#),
      2317 => to_slv(opcode_type, 16#09#),
      2318 => to_slv(opcode_type, 16#0C#),
      2319 => to_slv(opcode_type, 16#10#),
      2320 => to_slv(opcode_type, 16#06#),
      2321 => to_slv(opcode_type, 16#06#),
      2322 => to_slv(opcode_type, 16#08#),
      2323 => to_slv(opcode_type, 16#11#),
      2324 => to_slv(opcode_type, 16#10#),
      2325 => to_slv(opcode_type, 16#09#),
      2326 => to_slv(opcode_type, 16#0F#),
      2327 => to_slv(opcode_type, 16#0C#),
      2328 => to_slv(opcode_type, 16#07#),
      2329 => to_slv(opcode_type, 16#06#),
      2330 => to_slv(opcode_type, 16#8B#),
      2331 => to_slv(opcode_type, 16#0D#),
      2332 => to_slv(opcode_type, 16#08#),
      2333 => to_slv(opcode_type, 16#C8#),
      2334 => to_slv(opcode_type, 16#0F#),
      2335 to 2335 => (others => '0'),

      -- Program 73...
      2336 => to_slv(opcode_type, 16#08#),
      2337 => to_slv(opcode_type, 16#07#),
      2338 => to_slv(opcode_type, 16#07#),
      2339 => to_slv(opcode_type, 16#06#),
      2340 => to_slv(opcode_type, 16#0D#),
      2341 => to_slv(opcode_type, 16#0B#),
      2342 => to_slv(opcode_type, 16#09#),
      2343 => to_slv(opcode_type, 16#0B#),
      2344 => to_slv(opcode_type, 16#10#),
      2345 => to_slv(opcode_type, 16#08#),
      2346 => to_slv(opcode_type, 16#07#),
      2347 => to_slv(opcode_type, 16#0C#),
      2348 => to_slv(opcode_type, 16#0C#),
      2349 => to_slv(opcode_type, 16#07#),
      2350 => to_slv(opcode_type, 16#0F#),
      2351 => to_slv(opcode_type, 16#0B#),
      2352 => to_slv(opcode_type, 16#08#),
      2353 => to_slv(opcode_type, 16#09#),
      2354 => to_slv(opcode_type, 16#06#),
      2355 => to_slv(opcode_type, 16#10#),
      2356 => to_slv(opcode_type, 16#0C#),
      2357 => to_slv(opcode_type, 16#09#),
      2358 => to_slv(opcode_type, 16#11#),
      2359 => to_slv(opcode_type, 16#11#),
      2360 => to_slv(opcode_type, 16#07#),
      2361 => to_slv(opcode_type, 16#07#),
      2362 => to_slv(opcode_type, 16#0A#),
      2363 => to_slv(opcode_type, 16#11#),
      2364 => to_slv(opcode_type, 16#09#),
      2365 => to_slv(opcode_type, 16#0E#),
      2366 => to_slv(opcode_type, 16#0E#),
      2367 to 2367 => (others => '0'),

      -- Program 74...
      2368 => to_slv(opcode_type, 16#07#),
      2369 => to_slv(opcode_type, 16#09#),
      2370 => to_slv(opcode_type, 16#07#),
      2371 => to_slv(opcode_type, 16#08#),
      2372 => to_slv(opcode_type, 16#0C#),
      2373 => to_slv(opcode_type, 16#F8#),
      2374 => to_slv(opcode_type, 16#09#),
      2375 => to_slv(opcode_type, 16#11#),
      2376 => to_slv(opcode_type, 16#0D#),
      2377 => to_slv(opcode_type, 16#08#),
      2378 => to_slv(opcode_type, 16#08#),
      2379 => to_slv(opcode_type, 16#37#),
      2380 => to_slv(opcode_type, 16#0E#),
      2381 => to_slv(opcode_type, 16#07#),
      2382 => to_slv(opcode_type, 16#11#),
      2383 => to_slv(opcode_type, 16#0A#),
      2384 => to_slv(opcode_type, 16#07#),
      2385 => to_slv(opcode_type, 16#06#),
      2386 => to_slv(opcode_type, 16#06#),
      2387 => to_slv(opcode_type, 16#11#),
      2388 => to_slv(opcode_type, 16#E7#),
      2389 => to_slv(opcode_type, 16#09#),
      2390 => to_slv(opcode_type, 16#0A#),
      2391 => to_slv(opcode_type, 16#0C#),
      2392 => to_slv(opcode_type, 16#08#),
      2393 => to_slv(opcode_type, 16#08#),
      2394 => to_slv(opcode_type, 16#0C#),
      2395 => to_slv(opcode_type, 16#10#),
      2396 => to_slv(opcode_type, 16#08#),
      2397 => to_slv(opcode_type, 16#0C#),
      2398 => to_slv(opcode_type, 16#10#),
      2399 to 2399 => (others => '0'),

      -- Program 75...
      2400 => to_slv(opcode_type, 16#07#),
      2401 => to_slv(opcode_type, 16#06#),
      2402 => to_slv(opcode_type, 16#09#),
      2403 => to_slv(opcode_type, 16#07#),
      2404 => to_slv(opcode_type, 16#0A#),
      2405 => to_slv(opcode_type, 16#0A#),
      2406 => to_slv(opcode_type, 16#07#),
      2407 => to_slv(opcode_type, 16#11#),
      2408 => to_slv(opcode_type, 16#0F#),
      2409 => to_slv(opcode_type, 16#07#),
      2410 => to_slv(opcode_type, 16#09#),
      2411 => to_slv(opcode_type, 16#10#),
      2412 => to_slv(opcode_type, 16#11#),
      2413 => to_slv(opcode_type, 16#08#),
      2414 => to_slv(opcode_type, 16#0C#),
      2415 => to_slv(opcode_type, 16#11#),
      2416 => to_slv(opcode_type, 16#06#),
      2417 => to_slv(opcode_type, 16#06#),
      2418 => to_slv(opcode_type, 16#09#),
      2419 => to_slv(opcode_type, 16#0B#),
      2420 => to_slv(opcode_type, 16#0E#),
      2421 => to_slv(opcode_type, 16#09#),
      2422 => to_slv(opcode_type, 16#0D#),
      2423 => to_slv(opcode_type, 16#0F#),
      2424 => to_slv(opcode_type, 16#09#),
      2425 => to_slv(opcode_type, 16#06#),
      2426 => to_slv(opcode_type, 16#0C#),
      2427 => to_slv(opcode_type, 16#0D#),
      2428 => to_slv(opcode_type, 16#08#),
      2429 => to_slv(opcode_type, 16#0B#),
      2430 => to_slv(opcode_type, 16#11#),
      2431 to 2431 => (others => '0'),

      -- Program 76...
      2432 => to_slv(opcode_type, 16#06#),
      2433 => to_slv(opcode_type, 16#07#),
      2434 => to_slv(opcode_type, 16#08#),
      2435 => to_slv(opcode_type, 16#06#),
      2436 => to_slv(opcode_type, 16#0B#),
      2437 => to_slv(opcode_type, 16#37#),
      2438 => to_slv(opcode_type, 16#07#),
      2439 => to_slv(opcode_type, 16#11#),
      2440 => to_slv(opcode_type, 16#0D#),
      2441 => to_slv(opcode_type, 16#08#),
      2442 => to_slv(opcode_type, 16#08#),
      2443 => to_slv(opcode_type, 16#10#),
      2444 => to_slv(opcode_type, 16#0C#),
      2445 => to_slv(opcode_type, 16#06#),
      2446 => to_slv(opcode_type, 16#0F#),
      2447 => to_slv(opcode_type, 16#3A#),
      2448 => to_slv(opcode_type, 16#09#),
      2449 => to_slv(opcode_type, 16#08#),
      2450 => to_slv(opcode_type, 16#08#),
      2451 => to_slv(opcode_type, 16#0A#),
      2452 => to_slv(opcode_type, 16#0D#),
      2453 => to_slv(opcode_type, 16#08#),
      2454 => to_slv(opcode_type, 16#0B#),
      2455 => to_slv(opcode_type, 16#11#),
      2456 => to_slv(opcode_type, 16#07#),
      2457 => to_slv(opcode_type, 16#08#),
      2458 => to_slv(opcode_type, 16#0A#),
      2459 => to_slv(opcode_type, 16#0B#),
      2460 => to_slv(opcode_type, 16#08#),
      2461 => to_slv(opcode_type, 16#DA#),
      2462 => to_slv(opcode_type, 16#0A#),
      2463 to 2463 => (others => '0'),

      -- Program 77...
      2464 => to_slv(opcode_type, 16#06#),
      2465 => to_slv(opcode_type, 16#06#),
      2466 => to_slv(opcode_type, 16#09#),
      2467 => to_slv(opcode_type, 16#09#),
      2468 => to_slv(opcode_type, 16#10#),
      2469 => to_slv(opcode_type, 16#0D#),
      2470 => to_slv(opcode_type, 16#08#),
      2471 => to_slv(opcode_type, 16#10#),
      2472 => to_slv(opcode_type, 16#0B#),
      2473 => to_slv(opcode_type, 16#09#),
      2474 => to_slv(opcode_type, 16#06#),
      2475 => to_slv(opcode_type, 16#31#),
      2476 => to_slv(opcode_type, 16#0F#),
      2477 => to_slv(opcode_type, 16#07#),
      2478 => to_slv(opcode_type, 16#0E#),
      2479 => to_slv(opcode_type, 16#0C#),
      2480 => to_slv(opcode_type, 16#09#),
      2481 => to_slv(opcode_type, 16#06#),
      2482 => to_slv(opcode_type, 16#06#),
      2483 => to_slv(opcode_type, 16#11#),
      2484 => to_slv(opcode_type, 16#10#),
      2485 => to_slv(opcode_type, 16#07#),
      2486 => to_slv(opcode_type, 16#0F#),
      2487 => to_slv(opcode_type, 16#4E#),
      2488 => to_slv(opcode_type, 16#07#),
      2489 => to_slv(opcode_type, 16#08#),
      2490 => to_slv(opcode_type, 16#0E#),
      2491 => to_slv(opcode_type, 16#11#),
      2492 => to_slv(opcode_type, 16#07#),
      2493 => to_slv(opcode_type, 16#0E#),
      2494 => to_slv(opcode_type, 16#0D#),
      2495 to 2495 => (others => '0'),

      -- Program 78...
      2496 => to_slv(opcode_type, 16#09#),
      2497 => to_slv(opcode_type, 16#06#),
      2498 => to_slv(opcode_type, 16#07#),
      2499 => to_slv(opcode_type, 16#08#),
      2500 => to_slv(opcode_type, 16#0C#),
      2501 => to_slv(opcode_type, 16#0E#),
      2502 => to_slv(opcode_type, 16#07#),
      2503 => to_slv(opcode_type, 16#10#),
      2504 => to_slv(opcode_type, 16#0A#),
      2505 => to_slv(opcode_type, 16#06#),
      2506 => to_slv(opcode_type, 16#09#),
      2507 => to_slv(opcode_type, 16#0E#),
      2508 => to_slv(opcode_type, 16#0E#),
      2509 => to_slv(opcode_type, 16#06#),
      2510 => to_slv(opcode_type, 16#10#),
      2511 => to_slv(opcode_type, 16#10#),
      2512 => to_slv(opcode_type, 16#07#),
      2513 => to_slv(opcode_type, 16#06#),
      2514 => to_slv(opcode_type, 16#06#),
      2515 => to_slv(opcode_type, 16#10#),
      2516 => to_slv(opcode_type, 16#0A#),
      2517 => to_slv(opcode_type, 16#08#),
      2518 => to_slv(opcode_type, 16#0A#),
      2519 => to_slv(opcode_type, 16#0C#),
      2520 => to_slv(opcode_type, 16#07#),
      2521 => to_slv(opcode_type, 16#07#),
      2522 => to_slv(opcode_type, 16#0F#),
      2523 => to_slv(opcode_type, 16#1F#),
      2524 => to_slv(opcode_type, 16#06#),
      2525 => to_slv(opcode_type, 16#0E#),
      2526 => to_slv(opcode_type, 16#0A#),
      2527 to 2527 => (others => '0'),

      -- Program 79...
      2528 => to_slv(opcode_type, 16#06#),
      2529 => to_slv(opcode_type, 16#06#),
      2530 => to_slv(opcode_type, 16#06#),
      2531 => to_slv(opcode_type, 16#06#),
      2532 => to_slv(opcode_type, 16#0D#),
      2533 => to_slv(opcode_type, 16#B6#),
      2534 => to_slv(opcode_type, 16#06#),
      2535 => to_slv(opcode_type, 16#11#),
      2536 => to_slv(opcode_type, 16#0B#),
      2537 => to_slv(opcode_type, 16#07#),
      2538 => to_slv(opcode_type, 16#07#),
      2539 => to_slv(opcode_type, 16#D9#),
      2540 => to_slv(opcode_type, 16#0B#),
      2541 => to_slv(opcode_type, 16#06#),
      2542 => to_slv(opcode_type, 16#C5#),
      2543 => to_slv(opcode_type, 16#0A#),
      2544 => to_slv(opcode_type, 16#08#),
      2545 => to_slv(opcode_type, 16#09#),
      2546 => to_slv(opcode_type, 16#08#),
      2547 => to_slv(opcode_type, 16#10#),
      2548 => to_slv(opcode_type, 16#0D#),
      2549 => to_slv(opcode_type, 16#07#),
      2550 => to_slv(opcode_type, 16#65#),
      2551 => to_slv(opcode_type, 16#F8#),
      2552 => to_slv(opcode_type, 16#07#),
      2553 => to_slv(opcode_type, 16#08#),
      2554 => to_slv(opcode_type, 16#0E#),
      2555 => to_slv(opcode_type, 16#10#),
      2556 => to_slv(opcode_type, 16#08#),
      2557 => to_slv(opcode_type, 16#0E#),
      2558 => to_slv(opcode_type, 16#0A#),
      2559 to 2559 => (others => '0'),

      -- Program 80...
      2560 => to_slv(opcode_type, 16#06#),
      2561 => to_slv(opcode_type, 16#06#),
      2562 => to_slv(opcode_type, 16#07#),
      2563 => to_slv(opcode_type, 16#09#),
      2564 => to_slv(opcode_type, 16#0D#),
      2565 => to_slv(opcode_type, 16#7B#),
      2566 => to_slv(opcode_type, 16#08#),
      2567 => to_slv(opcode_type, 16#0F#),
      2568 => to_slv(opcode_type, 16#0E#),
      2569 => to_slv(opcode_type, 16#08#),
      2570 => to_slv(opcode_type, 16#08#),
      2571 => to_slv(opcode_type, 16#0D#),
      2572 => to_slv(opcode_type, 16#0C#),
      2573 => to_slv(opcode_type, 16#09#),
      2574 => to_slv(opcode_type, 16#11#),
      2575 => to_slv(opcode_type, 16#11#),
      2576 => to_slv(opcode_type, 16#08#),
      2577 => to_slv(opcode_type, 16#07#),
      2578 => to_slv(opcode_type, 16#08#),
      2579 => to_slv(opcode_type, 16#0E#),
      2580 => to_slv(opcode_type, 16#0E#),
      2581 => to_slv(opcode_type, 16#09#),
      2582 => to_slv(opcode_type, 16#0C#),
      2583 => to_slv(opcode_type, 16#0A#),
      2584 => to_slv(opcode_type, 16#07#),
      2585 => to_slv(opcode_type, 16#08#),
      2586 => to_slv(opcode_type, 16#0A#),
      2587 => to_slv(opcode_type, 16#10#),
      2588 => to_slv(opcode_type, 16#07#),
      2589 => to_slv(opcode_type, 16#0D#),
      2590 => to_slv(opcode_type, 16#0E#),
      2591 to 2591 => (others => '0'),

      -- Program 81...
      2592 => to_slv(opcode_type, 16#08#),
      2593 => to_slv(opcode_type, 16#06#),
      2594 => to_slv(opcode_type, 16#08#),
      2595 => to_slv(opcode_type, 16#06#),
      2596 => to_slv(opcode_type, 16#0A#),
      2597 => to_slv(opcode_type, 16#0A#),
      2598 => to_slv(opcode_type, 16#08#),
      2599 => to_slv(opcode_type, 16#0B#),
      2600 => to_slv(opcode_type, 16#0F#),
      2601 => to_slv(opcode_type, 16#06#),
      2602 => to_slv(opcode_type, 16#08#),
      2603 => to_slv(opcode_type, 16#0E#),
      2604 => to_slv(opcode_type, 16#0D#),
      2605 => to_slv(opcode_type, 16#07#),
      2606 => to_slv(opcode_type, 16#0E#),
      2607 => to_slv(opcode_type, 16#0D#),
      2608 => to_slv(opcode_type, 16#06#),
      2609 => to_slv(opcode_type, 16#07#),
      2610 => to_slv(opcode_type, 16#08#),
      2611 => to_slv(opcode_type, 16#0D#),
      2612 => to_slv(opcode_type, 16#0D#),
      2613 => to_slv(opcode_type, 16#06#),
      2614 => to_slv(opcode_type, 16#10#),
      2615 => to_slv(opcode_type, 16#0A#),
      2616 => to_slv(opcode_type, 16#09#),
      2617 => to_slv(opcode_type, 16#09#),
      2618 => to_slv(opcode_type, 16#0C#),
      2619 => to_slv(opcode_type, 16#11#),
      2620 => to_slv(opcode_type, 16#07#),
      2621 => to_slv(opcode_type, 16#0C#),
      2622 => to_slv(opcode_type, 16#0D#),
      2623 to 2623 => (others => '0'),

      -- Program 82...
      2624 => to_slv(opcode_type, 16#09#),
      2625 => to_slv(opcode_type, 16#06#),
      2626 => to_slv(opcode_type, 16#07#),
      2627 => to_slv(opcode_type, 16#07#),
      2628 => to_slv(opcode_type, 16#10#),
      2629 => to_slv(opcode_type, 16#0F#),
      2630 => to_slv(opcode_type, 16#06#),
      2631 => to_slv(opcode_type, 16#0F#),
      2632 => to_slv(opcode_type, 16#0F#),
      2633 => to_slv(opcode_type, 16#06#),
      2634 => to_slv(opcode_type, 16#08#),
      2635 => to_slv(opcode_type, 16#0A#),
      2636 => to_slv(opcode_type, 16#0D#),
      2637 => to_slv(opcode_type, 16#07#),
      2638 => to_slv(opcode_type, 16#0F#),
      2639 => to_slv(opcode_type, 16#0A#),
      2640 => to_slv(opcode_type, 16#09#),
      2641 => to_slv(opcode_type, 16#09#),
      2642 => to_slv(opcode_type, 16#09#),
      2643 => to_slv(opcode_type, 16#0A#),
      2644 => to_slv(opcode_type, 16#0D#),
      2645 => to_slv(opcode_type, 16#08#),
      2646 => to_slv(opcode_type, 16#0B#),
      2647 => to_slv(opcode_type, 16#E9#),
      2648 => to_slv(opcode_type, 16#09#),
      2649 => to_slv(opcode_type, 16#06#),
      2650 => to_slv(opcode_type, 16#10#),
      2651 => to_slv(opcode_type, 16#11#),
      2652 => to_slv(opcode_type, 16#08#),
      2653 => to_slv(opcode_type, 16#20#),
      2654 => to_slv(opcode_type, 16#0B#),
      2655 to 2655 => (others => '0'),

      -- Program 83...
      2656 => to_slv(opcode_type, 16#09#),
      2657 => to_slv(opcode_type, 16#09#),
      2658 => to_slv(opcode_type, 16#08#),
      2659 => to_slv(opcode_type, 16#07#),
      2660 => to_slv(opcode_type, 16#0B#),
      2661 => to_slv(opcode_type, 16#10#),
      2662 => to_slv(opcode_type, 16#06#),
      2663 => to_slv(opcode_type, 16#0F#),
      2664 => to_slv(opcode_type, 16#0A#),
      2665 => to_slv(opcode_type, 16#06#),
      2666 => to_slv(opcode_type, 16#07#),
      2667 => to_slv(opcode_type, 16#0B#),
      2668 => to_slv(opcode_type, 16#10#),
      2669 => to_slv(opcode_type, 16#08#),
      2670 => to_slv(opcode_type, 16#0D#),
      2671 => to_slv(opcode_type, 16#0C#),
      2672 => to_slv(opcode_type, 16#08#),
      2673 => to_slv(opcode_type, 16#08#),
      2674 => to_slv(opcode_type, 16#08#),
      2675 => to_slv(opcode_type, 16#11#),
      2676 => to_slv(opcode_type, 16#0A#),
      2677 => to_slv(opcode_type, 16#08#),
      2678 => to_slv(opcode_type, 16#10#),
      2679 => to_slv(opcode_type, 16#0D#),
      2680 => to_slv(opcode_type, 16#07#),
      2681 => to_slv(opcode_type, 16#09#),
      2682 => to_slv(opcode_type, 16#0D#),
      2683 => to_slv(opcode_type, 16#0F#),
      2684 => to_slv(opcode_type, 16#09#),
      2685 => to_slv(opcode_type, 16#0F#),
      2686 => to_slv(opcode_type, 16#0B#),
      2687 to 2687 => (others => '0'),

      -- Program 84...
      2688 => to_slv(opcode_type, 16#09#),
      2689 => to_slv(opcode_type, 16#08#),
      2690 => to_slv(opcode_type, 16#06#),
      2691 => to_slv(opcode_type, 16#07#),
      2692 => to_slv(opcode_type, 16#0B#),
      2693 => to_slv(opcode_type, 16#10#),
      2694 => to_slv(opcode_type, 16#08#),
      2695 => to_slv(opcode_type, 16#0F#),
      2696 => to_slv(opcode_type, 16#11#),
      2697 => to_slv(opcode_type, 16#07#),
      2698 => to_slv(opcode_type, 16#06#),
      2699 => to_slv(opcode_type, 16#0F#),
      2700 => to_slv(opcode_type, 16#EA#),
      2701 => to_slv(opcode_type, 16#08#),
      2702 => to_slv(opcode_type, 16#0D#),
      2703 => to_slv(opcode_type, 16#10#),
      2704 => to_slv(opcode_type, 16#06#),
      2705 => to_slv(opcode_type, 16#07#),
      2706 => to_slv(opcode_type, 16#07#),
      2707 => to_slv(opcode_type, 16#10#),
      2708 => to_slv(opcode_type, 16#11#),
      2709 => to_slv(opcode_type, 16#09#),
      2710 => to_slv(opcode_type, 16#0C#),
      2711 => to_slv(opcode_type, 16#10#),
      2712 => to_slv(opcode_type, 16#06#),
      2713 => to_slv(opcode_type, 16#08#),
      2714 => to_slv(opcode_type, 16#0B#),
      2715 => to_slv(opcode_type, 16#0B#),
      2716 => to_slv(opcode_type, 16#08#),
      2717 => to_slv(opcode_type, 16#53#),
      2718 => to_slv(opcode_type, 16#8F#),
      2719 to 2719 => (others => '0'),

      -- Program 85...
      2720 => to_slv(opcode_type, 16#06#),
      2721 => to_slv(opcode_type, 16#09#),
      2722 => to_slv(opcode_type, 16#09#),
      2723 => to_slv(opcode_type, 16#07#),
      2724 => to_slv(opcode_type, 16#0A#),
      2725 => to_slv(opcode_type, 16#0C#),
      2726 => to_slv(opcode_type, 16#07#),
      2727 => to_slv(opcode_type, 16#0D#),
      2728 => to_slv(opcode_type, 16#0B#),
      2729 => to_slv(opcode_type, 16#08#),
      2730 => to_slv(opcode_type, 16#08#),
      2731 => to_slv(opcode_type, 16#0B#),
      2732 => to_slv(opcode_type, 16#D1#),
      2733 => to_slv(opcode_type, 16#08#),
      2734 => to_slv(opcode_type, 16#0C#),
      2735 => to_slv(opcode_type, 16#0F#),
      2736 => to_slv(opcode_type, 16#08#),
      2737 => to_slv(opcode_type, 16#08#),
      2738 => to_slv(opcode_type, 16#06#),
      2739 => to_slv(opcode_type, 16#10#),
      2740 => to_slv(opcode_type, 16#0D#),
      2741 => to_slv(opcode_type, 16#07#),
      2742 => to_slv(opcode_type, 16#0F#),
      2743 => to_slv(opcode_type, 16#0F#),
      2744 => to_slv(opcode_type, 16#06#),
      2745 => to_slv(opcode_type, 16#08#),
      2746 => to_slv(opcode_type, 16#96#),
      2747 => to_slv(opcode_type, 16#0B#),
      2748 => to_slv(opcode_type, 16#08#),
      2749 => to_slv(opcode_type, 16#0D#),
      2750 => to_slv(opcode_type, 16#0D#),
      2751 to 2751 => (others => '0'),

      -- Program 86...
      2752 => to_slv(opcode_type, 16#07#),
      2753 => to_slv(opcode_type, 16#08#),
      2754 => to_slv(opcode_type, 16#06#),
      2755 => to_slv(opcode_type, 16#08#),
      2756 => to_slv(opcode_type, 16#52#),
      2757 => to_slv(opcode_type, 16#0B#),
      2758 => to_slv(opcode_type, 16#06#),
      2759 => to_slv(opcode_type, 16#0F#),
      2760 => to_slv(opcode_type, 16#0C#),
      2761 => to_slv(opcode_type, 16#06#),
      2762 => to_slv(opcode_type, 16#09#),
      2763 => to_slv(opcode_type, 16#0B#),
      2764 => to_slv(opcode_type, 16#0D#),
      2765 => to_slv(opcode_type, 16#09#),
      2766 => to_slv(opcode_type, 16#0C#),
      2767 => to_slv(opcode_type, 16#0A#),
      2768 => to_slv(opcode_type, 16#07#),
      2769 => to_slv(opcode_type, 16#09#),
      2770 => to_slv(opcode_type, 16#07#),
      2771 => to_slv(opcode_type, 16#0C#),
      2772 => to_slv(opcode_type, 16#0B#),
      2773 => to_slv(opcode_type, 16#07#),
      2774 => to_slv(opcode_type, 16#0A#),
      2775 => to_slv(opcode_type, 16#0C#),
      2776 => to_slv(opcode_type, 16#06#),
      2777 => to_slv(opcode_type, 16#07#),
      2778 => to_slv(opcode_type, 16#10#),
      2779 => to_slv(opcode_type, 16#0F#),
      2780 => to_slv(opcode_type, 16#09#),
      2781 => to_slv(opcode_type, 16#0E#),
      2782 => to_slv(opcode_type, 16#0F#),
      2783 to 2783 => (others => '0'),

      -- Program 87...
      2784 => to_slv(opcode_type, 16#09#),
      2785 => to_slv(opcode_type, 16#08#),
      2786 => to_slv(opcode_type, 16#07#),
      2787 => to_slv(opcode_type, 16#09#),
      2788 => to_slv(opcode_type, 16#0B#),
      2789 => to_slv(opcode_type, 16#0E#),
      2790 => to_slv(opcode_type, 16#06#),
      2791 => to_slv(opcode_type, 16#0E#),
      2792 => to_slv(opcode_type, 16#0E#),
      2793 => to_slv(opcode_type, 16#08#),
      2794 => to_slv(opcode_type, 16#07#),
      2795 => to_slv(opcode_type, 16#0F#),
      2796 => to_slv(opcode_type, 16#0B#),
      2797 => to_slv(opcode_type, 16#09#),
      2798 => to_slv(opcode_type, 16#0C#),
      2799 => to_slv(opcode_type, 16#0E#),
      2800 => to_slv(opcode_type, 16#06#),
      2801 => to_slv(opcode_type, 16#08#),
      2802 => to_slv(opcode_type, 16#06#),
      2803 => to_slv(opcode_type, 16#0F#),
      2804 => to_slv(opcode_type, 16#11#),
      2805 => to_slv(opcode_type, 16#09#),
      2806 => to_slv(opcode_type, 16#0E#),
      2807 => to_slv(opcode_type, 16#0E#),
      2808 => to_slv(opcode_type, 16#07#),
      2809 => to_slv(opcode_type, 16#09#),
      2810 => to_slv(opcode_type, 16#0D#),
      2811 => to_slv(opcode_type, 16#0F#),
      2812 => to_slv(opcode_type, 16#06#),
      2813 => to_slv(opcode_type, 16#0D#),
      2814 => to_slv(opcode_type, 16#0D#),
      2815 to 2815 => (others => '0'),

      -- Program 88...
      2816 => to_slv(opcode_type, 16#09#),
      2817 => to_slv(opcode_type, 16#09#),
      2818 => to_slv(opcode_type, 16#08#),
      2819 => to_slv(opcode_type, 16#09#),
      2820 => to_slv(opcode_type, 16#0E#),
      2821 => to_slv(opcode_type, 16#AE#),
      2822 => to_slv(opcode_type, 16#09#),
      2823 => to_slv(opcode_type, 16#0E#),
      2824 => to_slv(opcode_type, 16#10#),
      2825 => to_slv(opcode_type, 16#09#),
      2826 => to_slv(opcode_type, 16#08#),
      2827 => to_slv(opcode_type, 16#0A#),
      2828 => to_slv(opcode_type, 16#10#),
      2829 => to_slv(opcode_type, 16#06#),
      2830 => to_slv(opcode_type, 16#0D#),
      2831 => to_slv(opcode_type, 16#11#),
      2832 => to_slv(opcode_type, 16#07#),
      2833 => to_slv(opcode_type, 16#07#),
      2834 => to_slv(opcode_type, 16#09#),
      2835 => to_slv(opcode_type, 16#0E#),
      2836 => to_slv(opcode_type, 16#0C#),
      2837 => to_slv(opcode_type, 16#09#),
      2838 => to_slv(opcode_type, 16#0F#),
      2839 => to_slv(opcode_type, 16#10#),
      2840 => to_slv(opcode_type, 16#08#),
      2841 => to_slv(opcode_type, 16#07#),
      2842 => to_slv(opcode_type, 16#10#),
      2843 => to_slv(opcode_type, 16#0D#),
      2844 => to_slv(opcode_type, 16#08#),
      2845 => to_slv(opcode_type, 16#0B#),
      2846 => to_slv(opcode_type, 16#AC#),
      2847 to 2847 => (others => '0'),

      -- Program 89...
      2848 => to_slv(opcode_type, 16#09#),
      2849 => to_slv(opcode_type, 16#06#),
      2850 => to_slv(opcode_type, 16#06#),
      2851 => to_slv(opcode_type, 16#06#),
      2852 => to_slv(opcode_type, 16#0D#),
      2853 => to_slv(opcode_type, 16#0D#),
      2854 => to_slv(opcode_type, 16#09#),
      2855 => to_slv(opcode_type, 16#11#),
      2856 => to_slv(opcode_type, 16#11#),
      2857 => to_slv(opcode_type, 16#09#),
      2858 => to_slv(opcode_type, 16#06#),
      2859 => to_slv(opcode_type, 16#7D#),
      2860 => to_slv(opcode_type, 16#0C#),
      2861 => to_slv(opcode_type, 16#06#),
      2862 => to_slv(opcode_type, 16#0D#),
      2863 => to_slv(opcode_type, 16#0F#),
      2864 => to_slv(opcode_type, 16#08#),
      2865 => to_slv(opcode_type, 16#07#),
      2866 => to_slv(opcode_type, 16#08#),
      2867 => to_slv(opcode_type, 16#4A#),
      2868 => to_slv(opcode_type, 16#0E#),
      2869 => to_slv(opcode_type, 16#07#),
      2870 => to_slv(opcode_type, 16#0D#),
      2871 => to_slv(opcode_type, 16#0B#),
      2872 => to_slv(opcode_type, 16#07#),
      2873 => to_slv(opcode_type, 16#08#),
      2874 => to_slv(opcode_type, 16#0C#),
      2875 => to_slv(opcode_type, 16#0A#),
      2876 => to_slv(opcode_type, 16#06#),
      2877 => to_slv(opcode_type, 16#10#),
      2878 => to_slv(opcode_type, 16#0D#),
      2879 to 2879 => (others => '0'),

      -- Program 90...
      2880 => to_slv(opcode_type, 16#07#),
      2881 => to_slv(opcode_type, 16#08#),
      2882 => to_slv(opcode_type, 16#09#),
      2883 => to_slv(opcode_type, 16#06#),
      2884 => to_slv(opcode_type, 16#11#),
      2885 => to_slv(opcode_type, 16#0C#),
      2886 => to_slv(opcode_type, 16#07#),
      2887 => to_slv(opcode_type, 16#0B#),
      2888 => to_slv(opcode_type, 16#10#),
      2889 => to_slv(opcode_type, 16#07#),
      2890 => to_slv(opcode_type, 16#09#),
      2891 => to_slv(opcode_type, 16#0F#),
      2892 => to_slv(opcode_type, 16#0B#),
      2893 => to_slv(opcode_type, 16#06#),
      2894 => to_slv(opcode_type, 16#0F#),
      2895 => to_slv(opcode_type, 16#0D#),
      2896 => to_slv(opcode_type, 16#06#),
      2897 => to_slv(opcode_type, 16#07#),
      2898 => to_slv(opcode_type, 16#07#),
      2899 => to_slv(opcode_type, 16#0B#),
      2900 => to_slv(opcode_type, 16#10#),
      2901 => to_slv(opcode_type, 16#08#),
      2902 => to_slv(opcode_type, 16#10#),
      2903 => to_slv(opcode_type, 16#0E#),
      2904 => to_slv(opcode_type, 16#09#),
      2905 => to_slv(opcode_type, 16#08#),
      2906 => to_slv(opcode_type, 16#0F#),
      2907 => to_slv(opcode_type, 16#11#),
      2908 => to_slv(opcode_type, 16#06#),
      2909 => to_slv(opcode_type, 16#0E#),
      2910 => to_slv(opcode_type, 16#0A#),
      2911 to 2911 => (others => '0'),

      -- Program 91...
      2912 => to_slv(opcode_type, 16#09#),
      2913 => to_slv(opcode_type, 16#09#),
      2914 => to_slv(opcode_type, 16#06#),
      2915 => to_slv(opcode_type, 16#07#),
      2916 => to_slv(opcode_type, 16#0C#),
      2917 => to_slv(opcode_type, 16#0A#),
      2918 => to_slv(opcode_type, 16#08#),
      2919 => to_slv(opcode_type, 16#11#),
      2920 => to_slv(opcode_type, 16#0C#),
      2921 => to_slv(opcode_type, 16#06#),
      2922 => to_slv(opcode_type, 16#08#),
      2923 => to_slv(opcode_type, 16#0C#),
      2924 => to_slv(opcode_type, 16#0C#),
      2925 => to_slv(opcode_type, 16#08#),
      2926 => to_slv(opcode_type, 16#0F#),
      2927 => to_slv(opcode_type, 16#0B#),
      2928 => to_slv(opcode_type, 16#08#),
      2929 => to_slv(opcode_type, 16#06#),
      2930 => to_slv(opcode_type, 16#06#),
      2931 => to_slv(opcode_type, 16#0B#),
      2932 => to_slv(opcode_type, 16#10#),
      2933 => to_slv(opcode_type, 16#09#),
      2934 => to_slv(opcode_type, 16#0D#),
      2935 => to_slv(opcode_type, 16#11#),
      2936 => to_slv(opcode_type, 16#06#),
      2937 => to_slv(opcode_type, 16#08#),
      2938 => to_slv(opcode_type, 16#0E#),
      2939 => to_slv(opcode_type, 16#10#),
      2940 => to_slv(opcode_type, 16#08#),
      2941 => to_slv(opcode_type, 16#0D#),
      2942 => to_slv(opcode_type, 16#11#),
      2943 to 2943 => (others => '0'),

      -- Program 92...
      2944 => to_slv(opcode_type, 16#08#),
      2945 => to_slv(opcode_type, 16#08#),
      2946 => to_slv(opcode_type, 16#07#),
      2947 => to_slv(opcode_type, 16#07#),
      2948 => to_slv(opcode_type, 16#0F#),
      2949 => to_slv(opcode_type, 16#0F#),
      2950 => to_slv(opcode_type, 16#06#),
      2951 => to_slv(opcode_type, 16#0C#),
      2952 => to_slv(opcode_type, 16#11#),
      2953 => to_slv(opcode_type, 16#07#),
      2954 => to_slv(opcode_type, 16#08#),
      2955 => to_slv(opcode_type, 16#0B#),
      2956 => to_slv(opcode_type, 16#10#),
      2957 => to_slv(opcode_type, 16#06#),
      2958 => to_slv(opcode_type, 16#0C#),
      2959 => to_slv(opcode_type, 16#0E#),
      2960 => to_slv(opcode_type, 16#06#),
      2961 => to_slv(opcode_type, 16#06#),
      2962 => to_slv(opcode_type, 16#07#),
      2963 => to_slv(opcode_type, 16#0C#),
      2964 => to_slv(opcode_type, 16#0E#),
      2965 => to_slv(opcode_type, 16#06#),
      2966 => to_slv(opcode_type, 16#0B#),
      2967 => to_slv(opcode_type, 16#0A#),
      2968 => to_slv(opcode_type, 16#06#),
      2969 => to_slv(opcode_type, 16#09#),
      2970 => to_slv(opcode_type, 16#0D#),
      2971 => to_slv(opcode_type, 16#68#),
      2972 => to_slv(opcode_type, 16#06#),
      2973 => to_slv(opcode_type, 16#11#),
      2974 => to_slv(opcode_type, 16#0D#),
      2975 to 2975 => (others => '0'),

      -- Program 93...
      2976 => to_slv(opcode_type, 16#09#),
      2977 => to_slv(opcode_type, 16#09#),
      2978 => to_slv(opcode_type, 16#07#),
      2979 => to_slv(opcode_type, 16#09#),
      2980 => to_slv(opcode_type, 16#0F#),
      2981 => to_slv(opcode_type, 16#11#),
      2982 => to_slv(opcode_type, 16#06#),
      2983 => to_slv(opcode_type, 16#11#),
      2984 => to_slv(opcode_type, 16#0D#),
      2985 => to_slv(opcode_type, 16#06#),
      2986 => to_slv(opcode_type, 16#07#),
      2987 => to_slv(opcode_type, 16#0F#),
      2988 => to_slv(opcode_type, 16#0B#),
      2989 => to_slv(opcode_type, 16#08#),
      2990 => to_slv(opcode_type, 16#0C#),
      2991 => to_slv(opcode_type, 16#0A#),
      2992 => to_slv(opcode_type, 16#09#),
      2993 => to_slv(opcode_type, 16#07#),
      2994 => to_slv(opcode_type, 16#07#),
      2995 => to_slv(opcode_type, 16#10#),
      2996 => to_slv(opcode_type, 16#0B#),
      2997 => to_slv(opcode_type, 16#09#),
      2998 => to_slv(opcode_type, 16#0E#),
      2999 => to_slv(opcode_type, 16#89#),
      3000 => to_slv(opcode_type, 16#09#),
      3001 => to_slv(opcode_type, 16#09#),
      3002 => to_slv(opcode_type, 16#0A#),
      3003 => to_slv(opcode_type, 16#0A#),
      3004 => to_slv(opcode_type, 16#07#),
      3005 => to_slv(opcode_type, 16#10#),
      3006 => to_slv(opcode_type, 16#0E#),
      3007 to 3007 => (others => '0'),

      -- Program 94...
      3008 => to_slv(opcode_type, 16#07#),
      3009 => to_slv(opcode_type, 16#08#),
      3010 => to_slv(opcode_type, 16#06#),
      3011 => to_slv(opcode_type, 16#09#),
      3012 => to_slv(opcode_type, 16#0B#),
      3013 => to_slv(opcode_type, 16#0B#),
      3014 => to_slv(opcode_type, 16#08#),
      3015 => to_slv(opcode_type, 16#0A#),
      3016 => to_slv(opcode_type, 16#0C#),
      3017 => to_slv(opcode_type, 16#07#),
      3018 => to_slv(opcode_type, 16#08#),
      3019 => to_slv(opcode_type, 16#0E#),
      3020 => to_slv(opcode_type, 16#0F#),
      3021 => to_slv(opcode_type, 16#07#),
      3022 => to_slv(opcode_type, 16#B3#),
      3023 => to_slv(opcode_type, 16#11#),
      3024 => to_slv(opcode_type, 16#09#),
      3025 => to_slv(opcode_type, 16#08#),
      3026 => to_slv(opcode_type, 16#09#),
      3027 => to_slv(opcode_type, 16#0D#),
      3028 => to_slv(opcode_type, 16#0C#),
      3029 => to_slv(opcode_type, 16#07#),
      3030 => to_slv(opcode_type, 16#0F#),
      3031 => to_slv(opcode_type, 16#10#),
      3032 => to_slv(opcode_type, 16#09#),
      3033 => to_slv(opcode_type, 16#08#),
      3034 => to_slv(opcode_type, 16#0A#),
      3035 => to_slv(opcode_type, 16#0D#),
      3036 => to_slv(opcode_type, 16#06#),
      3037 => to_slv(opcode_type, 16#0B#),
      3038 => to_slv(opcode_type, 16#0B#),
      3039 to 3039 => (others => '0'),

      -- Program 95...
      3040 => to_slv(opcode_type, 16#07#),
      3041 => to_slv(opcode_type, 16#06#),
      3042 => to_slv(opcode_type, 16#09#),
      3043 => to_slv(opcode_type, 16#07#),
      3044 => to_slv(opcode_type, 16#0B#),
      3045 => to_slv(opcode_type, 16#0D#),
      3046 => to_slv(opcode_type, 16#07#),
      3047 => to_slv(opcode_type, 16#AC#),
      3048 => to_slv(opcode_type, 16#0F#),
      3049 => to_slv(opcode_type, 16#06#),
      3050 => to_slv(opcode_type, 16#08#),
      3051 => to_slv(opcode_type, 16#0C#),
      3052 => to_slv(opcode_type, 16#0F#),
      3053 => to_slv(opcode_type, 16#09#),
      3054 => to_slv(opcode_type, 16#10#),
      3055 => to_slv(opcode_type, 16#0B#),
      3056 => to_slv(opcode_type, 16#08#),
      3057 => to_slv(opcode_type, 16#06#),
      3058 => to_slv(opcode_type, 16#06#),
      3059 => to_slv(opcode_type, 16#11#),
      3060 => to_slv(opcode_type, 16#10#),
      3061 => to_slv(opcode_type, 16#06#),
      3062 => to_slv(opcode_type, 16#0B#),
      3063 => to_slv(opcode_type, 16#0F#),
      3064 => to_slv(opcode_type, 16#09#),
      3065 => to_slv(opcode_type, 16#06#),
      3066 => to_slv(opcode_type, 16#11#),
      3067 => to_slv(opcode_type, 16#0B#),
      3068 => to_slv(opcode_type, 16#09#),
      3069 => to_slv(opcode_type, 16#10#),
      3070 => to_slv(opcode_type, 16#0B#),
      3071 to 3071 => (others => '0'),

      -- Program 96...
      3072 => to_slv(opcode_type, 16#07#),
      3073 => to_slv(opcode_type, 16#08#),
      3074 => to_slv(opcode_type, 16#09#),
      3075 => to_slv(opcode_type, 16#09#),
      3076 => to_slv(opcode_type, 16#79#),
      3077 => to_slv(opcode_type, 16#0A#),
      3078 => to_slv(opcode_type, 16#06#),
      3079 => to_slv(opcode_type, 16#0C#),
      3080 => to_slv(opcode_type, 16#0F#),
      3081 => to_slv(opcode_type, 16#07#),
      3082 => to_slv(opcode_type, 16#09#),
      3083 => to_slv(opcode_type, 16#0A#),
      3084 => to_slv(opcode_type, 16#0F#),
      3085 => to_slv(opcode_type, 16#08#),
      3086 => to_slv(opcode_type, 16#0A#),
      3087 => to_slv(opcode_type, 16#0E#),
      3088 => to_slv(opcode_type, 16#09#),
      3089 => to_slv(opcode_type, 16#09#),
      3090 => to_slv(opcode_type, 16#07#),
      3091 => to_slv(opcode_type, 16#0A#),
      3092 => to_slv(opcode_type, 16#10#),
      3093 => to_slv(opcode_type, 16#08#),
      3094 => to_slv(opcode_type, 16#10#),
      3095 => to_slv(opcode_type, 16#0B#),
      3096 => to_slv(opcode_type, 16#09#),
      3097 => to_slv(opcode_type, 16#06#),
      3098 => to_slv(opcode_type, 16#0C#),
      3099 => to_slv(opcode_type, 16#11#),
      3100 => to_slv(opcode_type, 16#08#),
      3101 => to_slv(opcode_type, 16#11#),
      3102 => to_slv(opcode_type, 16#0E#),
      3103 to 3103 => (others => '0'),

      -- Program 97...
      3104 => to_slv(opcode_type, 16#06#),
      3105 => to_slv(opcode_type, 16#06#),
      3106 => to_slv(opcode_type, 16#08#),
      3107 => to_slv(opcode_type, 16#09#),
      3108 => to_slv(opcode_type, 16#0E#),
      3109 => to_slv(opcode_type, 16#0B#),
      3110 => to_slv(opcode_type, 16#09#),
      3111 => to_slv(opcode_type, 16#0B#),
      3112 => to_slv(opcode_type, 16#11#),
      3113 => to_slv(opcode_type, 16#06#),
      3114 => to_slv(opcode_type, 16#06#),
      3115 => to_slv(opcode_type, 16#0D#),
      3116 => to_slv(opcode_type, 16#0C#),
      3117 => to_slv(opcode_type, 16#08#),
      3118 => to_slv(opcode_type, 16#10#),
      3119 => to_slv(opcode_type, 16#10#),
      3120 => to_slv(opcode_type, 16#08#),
      3121 => to_slv(opcode_type, 16#06#),
      3122 => to_slv(opcode_type, 16#08#),
      3123 => to_slv(opcode_type, 16#11#),
      3124 => to_slv(opcode_type, 16#0F#),
      3125 => to_slv(opcode_type, 16#06#),
      3126 => to_slv(opcode_type, 16#0C#),
      3127 => to_slv(opcode_type, 16#0F#),
      3128 => to_slv(opcode_type, 16#09#),
      3129 => to_slv(opcode_type, 16#08#),
      3130 => to_slv(opcode_type, 16#0A#),
      3131 => to_slv(opcode_type, 16#0C#),
      3132 => to_slv(opcode_type, 16#09#),
      3133 => to_slv(opcode_type, 16#0C#),
      3134 => to_slv(opcode_type, 16#0B#),
      3135 to 3135 => (others => '0'),

      -- Program 98...
      3136 => to_slv(opcode_type, 16#07#),
      3137 => to_slv(opcode_type, 16#07#),
      3138 => to_slv(opcode_type, 16#08#),
      3139 => to_slv(opcode_type, 16#09#),
      3140 => to_slv(opcode_type, 16#11#),
      3141 => to_slv(opcode_type, 16#11#),
      3142 => to_slv(opcode_type, 16#08#),
      3143 => to_slv(opcode_type, 16#11#),
      3144 => to_slv(opcode_type, 16#10#),
      3145 => to_slv(opcode_type, 16#09#),
      3146 => to_slv(opcode_type, 16#09#),
      3147 => to_slv(opcode_type, 16#0A#),
      3148 => to_slv(opcode_type, 16#E8#),
      3149 => to_slv(opcode_type, 16#08#),
      3150 => to_slv(opcode_type, 16#0A#),
      3151 => to_slv(opcode_type, 16#9D#),
      3152 => to_slv(opcode_type, 16#06#),
      3153 => to_slv(opcode_type, 16#07#),
      3154 => to_slv(opcode_type, 16#08#),
      3155 => to_slv(opcode_type, 16#0D#),
      3156 => to_slv(opcode_type, 16#0C#),
      3157 => to_slv(opcode_type, 16#09#),
      3158 => to_slv(opcode_type, 16#0E#),
      3159 => to_slv(opcode_type, 16#0C#),
      3160 => to_slv(opcode_type, 16#07#),
      3161 => to_slv(opcode_type, 16#06#),
      3162 => to_slv(opcode_type, 16#10#),
      3163 => to_slv(opcode_type, 16#0A#),
      3164 => to_slv(opcode_type, 16#06#),
      3165 => to_slv(opcode_type, 16#AC#),
      3166 => to_slv(opcode_type, 16#11#),
      3167 to 3167 => (others => '0'),

      -- Program 99...
      3168 => to_slv(opcode_type, 16#09#),
      3169 => to_slv(opcode_type, 16#06#),
      3170 => to_slv(opcode_type, 16#08#),
      3171 => to_slv(opcode_type, 16#09#),
      3172 => to_slv(opcode_type, 16#0B#),
      3173 => to_slv(opcode_type, 16#0B#),
      3174 => to_slv(opcode_type, 16#08#),
      3175 => to_slv(opcode_type, 16#FE#),
      3176 => to_slv(opcode_type, 16#0C#),
      3177 => to_slv(opcode_type, 16#06#),
      3178 => to_slv(opcode_type, 16#07#),
      3179 => to_slv(opcode_type, 16#11#),
      3180 => to_slv(opcode_type, 16#0F#),
      3181 => to_slv(opcode_type, 16#07#),
      3182 => to_slv(opcode_type, 16#0B#),
      3183 => to_slv(opcode_type, 16#0F#),
      3184 => to_slv(opcode_type, 16#06#),
      3185 => to_slv(opcode_type, 16#06#),
      3186 => to_slv(opcode_type, 16#09#),
      3187 => to_slv(opcode_type, 16#0E#),
      3188 => to_slv(opcode_type, 16#11#),
      3189 => to_slv(opcode_type, 16#08#),
      3190 => to_slv(opcode_type, 16#0C#),
      3191 => to_slv(opcode_type, 16#0D#),
      3192 => to_slv(opcode_type, 16#07#),
      3193 => to_slv(opcode_type, 16#07#),
      3194 => to_slv(opcode_type, 16#0B#),
      3195 => to_slv(opcode_type, 16#0E#),
      3196 => to_slv(opcode_type, 16#09#),
      3197 => to_slv(opcode_type, 16#10#),
      3198 => to_slv(opcode_type, 16#10#),
      3199 to 3199 => (others => '0'),

      -- Program 100...
      3200 => to_slv(opcode_type, 16#09#),
      3201 => to_slv(opcode_type, 16#08#),
      3202 => to_slv(opcode_type, 16#09#),
      3203 => to_slv(opcode_type, 16#09#),
      3204 => to_slv(opcode_type, 16#C7#),
      3205 => to_slv(opcode_type, 16#0F#),
      3206 => to_slv(opcode_type, 16#09#),
      3207 => to_slv(opcode_type, 16#CC#),
      3208 => to_slv(opcode_type, 16#0E#),
      3209 => to_slv(opcode_type, 16#06#),
      3210 => to_slv(opcode_type, 16#08#),
      3211 => to_slv(opcode_type, 16#0D#),
      3212 => to_slv(opcode_type, 16#FB#),
      3213 => to_slv(opcode_type, 16#06#),
      3214 => to_slv(opcode_type, 16#0D#),
      3215 => to_slv(opcode_type, 16#0F#),
      3216 => to_slv(opcode_type, 16#06#),
      3217 => to_slv(opcode_type, 16#09#),
      3218 => to_slv(opcode_type, 16#07#),
      3219 => to_slv(opcode_type, 16#0C#),
      3220 => to_slv(opcode_type, 16#0C#),
      3221 => to_slv(opcode_type, 16#08#),
      3222 => to_slv(opcode_type, 16#11#),
      3223 => to_slv(opcode_type, 16#11#),
      3224 => to_slv(opcode_type, 16#09#),
      3225 => to_slv(opcode_type, 16#06#),
      3226 => to_slv(opcode_type, 16#11#),
      3227 => to_slv(opcode_type, 16#0E#),
      3228 => to_slv(opcode_type, 16#09#),
      3229 => to_slv(opcode_type, 16#0C#),
      3230 => to_slv(opcode_type, 16#0F#),
      3231 to 3231 => (others => '0'),

      -- Program 101...
      3232 => to_slv(opcode_type, 16#07#),
      3233 => to_slv(opcode_type, 16#09#),
      3234 => to_slv(opcode_type, 16#07#),
      3235 => to_slv(opcode_type, 16#07#),
      3236 => to_slv(opcode_type, 16#11#),
      3237 => to_slv(opcode_type, 16#0F#),
      3238 => to_slv(opcode_type, 16#08#),
      3239 => to_slv(opcode_type, 16#10#),
      3240 => to_slv(opcode_type, 16#0B#),
      3241 => to_slv(opcode_type, 16#09#),
      3242 => to_slv(opcode_type, 16#06#),
      3243 => to_slv(opcode_type, 16#0F#),
      3244 => to_slv(opcode_type, 16#0C#),
      3245 => to_slv(opcode_type, 16#09#),
      3246 => to_slv(opcode_type, 16#11#),
      3247 => to_slv(opcode_type, 16#10#),
      3248 => to_slv(opcode_type, 16#09#),
      3249 => to_slv(opcode_type, 16#09#),
      3250 => to_slv(opcode_type, 16#08#),
      3251 => to_slv(opcode_type, 16#0E#),
      3252 => to_slv(opcode_type, 16#0B#),
      3253 => to_slv(opcode_type, 16#09#),
      3254 => to_slv(opcode_type, 16#0E#),
      3255 => to_slv(opcode_type, 16#0A#),
      3256 => to_slv(opcode_type, 16#08#),
      3257 => to_slv(opcode_type, 16#08#),
      3258 => to_slv(opcode_type, 16#0C#),
      3259 => to_slv(opcode_type, 16#11#),
      3260 => to_slv(opcode_type, 16#09#),
      3261 => to_slv(opcode_type, 16#11#),
      3262 => to_slv(opcode_type, 16#D2#),
      3263 to 3263 => (others => '0'),

      -- Program 102...
      3264 => to_slv(opcode_type, 16#09#),
      3265 => to_slv(opcode_type, 16#07#),
      3266 => to_slv(opcode_type, 16#09#),
      3267 => to_slv(opcode_type, 16#07#),
      3268 => to_slv(opcode_type, 16#0A#),
      3269 => to_slv(opcode_type, 16#11#),
      3270 => to_slv(opcode_type, 16#07#),
      3271 => to_slv(opcode_type, 16#0D#),
      3272 => to_slv(opcode_type, 16#5E#),
      3273 => to_slv(opcode_type, 16#07#),
      3274 => to_slv(opcode_type, 16#06#),
      3275 => to_slv(opcode_type, 16#0F#),
      3276 => to_slv(opcode_type, 16#0C#),
      3277 => to_slv(opcode_type, 16#09#),
      3278 => to_slv(opcode_type, 16#0C#),
      3279 => to_slv(opcode_type, 16#0F#),
      3280 => to_slv(opcode_type, 16#09#),
      3281 => to_slv(opcode_type, 16#08#),
      3282 => to_slv(opcode_type, 16#08#),
      3283 => to_slv(opcode_type, 16#0C#),
      3284 => to_slv(opcode_type, 16#11#),
      3285 => to_slv(opcode_type, 16#08#),
      3286 => to_slv(opcode_type, 16#0E#),
      3287 => to_slv(opcode_type, 16#5D#),
      3288 => to_slv(opcode_type, 16#08#),
      3289 => to_slv(opcode_type, 16#06#),
      3290 => to_slv(opcode_type, 16#0D#),
      3291 => to_slv(opcode_type, 16#0D#),
      3292 => to_slv(opcode_type, 16#06#),
      3293 => to_slv(opcode_type, 16#36#),
      3294 => to_slv(opcode_type, 16#0A#),
      3295 to 3295 => (others => '0'),

      -- Program 103...
      3296 => to_slv(opcode_type, 16#08#),
      3297 => to_slv(opcode_type, 16#08#),
      3298 => to_slv(opcode_type, 16#07#),
      3299 => to_slv(opcode_type, 16#07#),
      3300 => to_slv(opcode_type, 16#0F#),
      3301 => to_slv(opcode_type, 16#B7#),
      3302 => to_slv(opcode_type, 16#07#),
      3303 => to_slv(opcode_type, 16#11#),
      3304 => to_slv(opcode_type, 16#E2#),
      3305 => to_slv(opcode_type, 16#06#),
      3306 => to_slv(opcode_type, 16#08#),
      3307 => to_slv(opcode_type, 16#10#),
      3308 => to_slv(opcode_type, 16#0C#),
      3309 => to_slv(opcode_type, 16#08#),
      3310 => to_slv(opcode_type, 16#0D#),
      3311 => to_slv(opcode_type, 16#0A#),
      3312 => to_slv(opcode_type, 16#06#),
      3313 => to_slv(opcode_type, 16#06#),
      3314 => to_slv(opcode_type, 16#08#),
      3315 => to_slv(opcode_type, 16#10#),
      3316 => to_slv(opcode_type, 16#11#),
      3317 => to_slv(opcode_type, 16#06#),
      3318 => to_slv(opcode_type, 16#0B#),
      3319 => to_slv(opcode_type, 16#0C#),
      3320 => to_slv(opcode_type, 16#09#),
      3321 => to_slv(opcode_type, 16#09#),
      3322 => to_slv(opcode_type, 16#0B#),
      3323 => to_slv(opcode_type, 16#FE#),
      3324 => to_slv(opcode_type, 16#08#),
      3325 => to_slv(opcode_type, 16#0E#),
      3326 => to_slv(opcode_type, 16#0A#),
      3327 to 3327 => (others => '0'),

      -- Program 104...
      3328 => to_slv(opcode_type, 16#06#),
      3329 => to_slv(opcode_type, 16#09#),
      3330 => to_slv(opcode_type, 16#08#),
      3331 => to_slv(opcode_type, 16#08#),
      3332 => to_slv(opcode_type, 16#0A#),
      3333 => to_slv(opcode_type, 16#0D#),
      3334 => to_slv(opcode_type, 16#06#),
      3335 => to_slv(opcode_type, 16#0D#),
      3336 => to_slv(opcode_type, 16#0B#),
      3337 => to_slv(opcode_type, 16#09#),
      3338 => to_slv(opcode_type, 16#09#),
      3339 => to_slv(opcode_type, 16#0F#),
      3340 => to_slv(opcode_type, 16#0F#),
      3341 => to_slv(opcode_type, 16#07#),
      3342 => to_slv(opcode_type, 16#0A#),
      3343 => to_slv(opcode_type, 16#0F#),
      3344 => to_slv(opcode_type, 16#06#),
      3345 => to_slv(opcode_type, 16#08#),
      3346 => to_slv(opcode_type, 16#07#),
      3347 => to_slv(opcode_type, 16#0E#),
      3348 => to_slv(opcode_type, 16#10#),
      3349 => to_slv(opcode_type, 16#06#),
      3350 => to_slv(opcode_type, 16#0C#),
      3351 => to_slv(opcode_type, 16#11#),
      3352 => to_slv(opcode_type, 16#09#),
      3353 => to_slv(opcode_type, 16#07#),
      3354 => to_slv(opcode_type, 16#0A#),
      3355 => to_slv(opcode_type, 16#10#),
      3356 => to_slv(opcode_type, 16#06#),
      3357 => to_slv(opcode_type, 16#0D#),
      3358 => to_slv(opcode_type, 16#0A#),
      3359 to 3359 => (others => '0'),

      -- Program 105...
      3360 => to_slv(opcode_type, 16#08#),
      3361 => to_slv(opcode_type, 16#08#),
      3362 => to_slv(opcode_type, 16#06#),
      3363 => to_slv(opcode_type, 16#07#),
      3364 => to_slv(opcode_type, 16#D9#),
      3365 => to_slv(opcode_type, 16#0E#),
      3366 => to_slv(opcode_type, 16#07#),
      3367 => to_slv(opcode_type, 16#10#),
      3368 => to_slv(opcode_type, 16#11#),
      3369 => to_slv(opcode_type, 16#07#),
      3370 => to_slv(opcode_type, 16#08#),
      3371 => to_slv(opcode_type, 16#0B#),
      3372 => to_slv(opcode_type, 16#0C#),
      3373 => to_slv(opcode_type, 16#09#),
      3374 => to_slv(opcode_type, 16#11#),
      3375 => to_slv(opcode_type, 16#10#),
      3376 => to_slv(opcode_type, 16#08#),
      3377 => to_slv(opcode_type, 16#09#),
      3378 => to_slv(opcode_type, 16#07#),
      3379 => to_slv(opcode_type, 16#0E#),
      3380 => to_slv(opcode_type, 16#0F#),
      3381 => to_slv(opcode_type, 16#08#),
      3382 => to_slv(opcode_type, 16#0C#),
      3383 => to_slv(opcode_type, 16#DD#),
      3384 => to_slv(opcode_type, 16#06#),
      3385 => to_slv(opcode_type, 16#09#),
      3386 => to_slv(opcode_type, 16#0D#),
      3387 => to_slv(opcode_type, 16#0D#),
      3388 => to_slv(opcode_type, 16#08#),
      3389 => to_slv(opcode_type, 16#11#),
      3390 => to_slv(opcode_type, 16#0D#),
      3391 to 3391 => (others => '0'),

      -- Program 106...
      3392 => to_slv(opcode_type, 16#07#),
      3393 => to_slv(opcode_type, 16#08#),
      3394 => to_slv(opcode_type, 16#07#),
      3395 => to_slv(opcode_type, 16#09#),
      3396 => to_slv(opcode_type, 16#10#),
      3397 => to_slv(opcode_type, 16#0C#),
      3398 => to_slv(opcode_type, 16#07#),
      3399 => to_slv(opcode_type, 16#0A#),
      3400 => to_slv(opcode_type, 16#10#),
      3401 => to_slv(opcode_type, 16#06#),
      3402 => to_slv(opcode_type, 16#08#),
      3403 => to_slv(opcode_type, 16#0F#),
      3404 => to_slv(opcode_type, 16#0B#),
      3405 => to_slv(opcode_type, 16#07#),
      3406 => to_slv(opcode_type, 16#0A#),
      3407 => to_slv(opcode_type, 16#11#),
      3408 => to_slv(opcode_type, 16#08#),
      3409 => to_slv(opcode_type, 16#09#),
      3410 => to_slv(opcode_type, 16#06#),
      3411 => to_slv(opcode_type, 16#10#),
      3412 => to_slv(opcode_type, 16#0C#),
      3413 => to_slv(opcode_type, 16#09#),
      3414 => to_slv(opcode_type, 16#0E#),
      3415 => to_slv(opcode_type, 16#10#),
      3416 => to_slv(opcode_type, 16#09#),
      3417 => to_slv(opcode_type, 16#06#),
      3418 => to_slv(opcode_type, 16#0B#),
      3419 => to_slv(opcode_type, 16#0C#),
      3420 => to_slv(opcode_type, 16#06#),
      3421 => to_slv(opcode_type, 16#10#),
      3422 => to_slv(opcode_type, 16#0C#),
      3423 to 3423 => (others => '0'),

      -- Program 107...
      3424 => to_slv(opcode_type, 16#07#),
      3425 => to_slv(opcode_type, 16#08#),
      3426 => to_slv(opcode_type, 16#09#),
      3427 => to_slv(opcode_type, 16#08#),
      3428 => to_slv(opcode_type, 16#0B#),
      3429 => to_slv(opcode_type, 16#10#),
      3430 => to_slv(opcode_type, 16#09#),
      3431 => to_slv(opcode_type, 16#EC#),
      3432 => to_slv(opcode_type, 16#11#),
      3433 => to_slv(opcode_type, 16#09#),
      3434 => to_slv(opcode_type, 16#08#),
      3435 => to_slv(opcode_type, 16#0F#),
      3436 => to_slv(opcode_type, 16#0B#),
      3437 => to_slv(opcode_type, 16#07#),
      3438 => to_slv(opcode_type, 16#0C#),
      3439 => to_slv(opcode_type, 16#21#),
      3440 => to_slv(opcode_type, 16#09#),
      3441 => to_slv(opcode_type, 16#09#),
      3442 => to_slv(opcode_type, 16#07#),
      3443 => to_slv(opcode_type, 16#0B#),
      3444 => to_slv(opcode_type, 16#0A#),
      3445 => to_slv(opcode_type, 16#08#),
      3446 => to_slv(opcode_type, 16#10#),
      3447 => to_slv(opcode_type, 16#0C#),
      3448 => to_slv(opcode_type, 16#07#),
      3449 => to_slv(opcode_type, 16#07#),
      3450 => to_slv(opcode_type, 16#29#),
      3451 => to_slv(opcode_type, 16#0B#),
      3452 => to_slv(opcode_type, 16#09#),
      3453 => to_slv(opcode_type, 16#11#),
      3454 => to_slv(opcode_type, 16#0D#),
      3455 to 3455 => (others => '0'),

      -- Program 108...
      3456 => to_slv(opcode_type, 16#06#),
      3457 => to_slv(opcode_type, 16#09#),
      3458 => to_slv(opcode_type, 16#06#),
      3459 => to_slv(opcode_type, 16#08#),
      3460 => to_slv(opcode_type, 16#0E#),
      3461 => to_slv(opcode_type, 16#0C#),
      3462 => to_slv(opcode_type, 16#09#),
      3463 => to_slv(opcode_type, 16#11#),
      3464 => to_slv(opcode_type, 16#0A#),
      3465 => to_slv(opcode_type, 16#09#),
      3466 => to_slv(opcode_type, 16#09#),
      3467 => to_slv(opcode_type, 16#0B#),
      3468 => to_slv(opcode_type, 16#0B#),
      3469 => to_slv(opcode_type, 16#09#),
      3470 => to_slv(opcode_type, 16#0A#),
      3471 => to_slv(opcode_type, 16#0F#),
      3472 => to_slv(opcode_type, 16#07#),
      3473 => to_slv(opcode_type, 16#09#),
      3474 => to_slv(opcode_type, 16#08#),
      3475 => to_slv(opcode_type, 16#0A#),
      3476 => to_slv(opcode_type, 16#0E#),
      3477 => to_slv(opcode_type, 16#08#),
      3478 => to_slv(opcode_type, 16#0E#),
      3479 => to_slv(opcode_type, 16#0E#),
      3480 => to_slv(opcode_type, 16#09#),
      3481 => to_slv(opcode_type, 16#08#),
      3482 => to_slv(opcode_type, 16#0A#),
      3483 => to_slv(opcode_type, 16#17#),
      3484 => to_slv(opcode_type, 16#07#),
      3485 => to_slv(opcode_type, 16#0B#),
      3486 => to_slv(opcode_type, 16#86#),
      3487 to 3487 => (others => '0'),

      -- Program 109...
      3488 => to_slv(opcode_type, 16#07#),
      3489 => to_slv(opcode_type, 16#09#),
      3490 => to_slv(opcode_type, 16#08#),
      3491 => to_slv(opcode_type, 16#06#),
      3492 => to_slv(opcode_type, 16#0E#),
      3493 => to_slv(opcode_type, 16#11#),
      3494 => to_slv(opcode_type, 16#08#),
      3495 => to_slv(opcode_type, 16#0C#),
      3496 => to_slv(opcode_type, 16#9B#),
      3497 => to_slv(opcode_type, 16#09#),
      3498 => to_slv(opcode_type, 16#08#),
      3499 => to_slv(opcode_type, 16#0C#),
      3500 => to_slv(opcode_type, 16#0F#),
      3501 => to_slv(opcode_type, 16#07#),
      3502 => to_slv(opcode_type, 16#24#),
      3503 => to_slv(opcode_type, 16#0D#),
      3504 => to_slv(opcode_type, 16#06#),
      3505 => to_slv(opcode_type, 16#09#),
      3506 => to_slv(opcode_type, 16#07#),
      3507 => to_slv(opcode_type, 16#0B#),
      3508 => to_slv(opcode_type, 16#0A#),
      3509 => to_slv(opcode_type, 16#06#),
      3510 => to_slv(opcode_type, 16#47#),
      3511 => to_slv(opcode_type, 16#10#),
      3512 => to_slv(opcode_type, 16#07#),
      3513 => to_slv(opcode_type, 16#08#),
      3514 => to_slv(opcode_type, 16#11#),
      3515 => to_slv(opcode_type, 16#0B#),
      3516 => to_slv(opcode_type, 16#08#),
      3517 => to_slv(opcode_type, 16#0E#),
      3518 => to_slv(opcode_type, 16#10#),
      3519 to 3519 => (others => '0'),

      -- Program 110...
      3520 => to_slv(opcode_type, 16#07#),
      3521 => to_slv(opcode_type, 16#06#),
      3522 => to_slv(opcode_type, 16#09#),
      3523 => to_slv(opcode_type, 16#07#),
      3524 => to_slv(opcode_type, 16#11#),
      3525 => to_slv(opcode_type, 16#10#),
      3526 => to_slv(opcode_type, 16#06#),
      3527 => to_slv(opcode_type, 16#0E#),
      3528 => to_slv(opcode_type, 16#0A#),
      3529 => to_slv(opcode_type, 16#06#),
      3530 => to_slv(opcode_type, 16#08#),
      3531 => to_slv(opcode_type, 16#0A#),
      3532 => to_slv(opcode_type, 16#10#),
      3533 => to_slv(opcode_type, 16#08#),
      3534 => to_slv(opcode_type, 16#10#),
      3535 => to_slv(opcode_type, 16#10#),
      3536 => to_slv(opcode_type, 16#08#),
      3537 => to_slv(opcode_type, 16#09#),
      3538 => to_slv(opcode_type, 16#08#),
      3539 => to_slv(opcode_type, 16#0B#),
      3540 => to_slv(opcode_type, 16#0F#),
      3541 => to_slv(opcode_type, 16#09#),
      3542 => to_slv(opcode_type, 16#0E#),
      3543 => to_slv(opcode_type, 16#B1#),
      3544 => to_slv(opcode_type, 16#06#),
      3545 => to_slv(opcode_type, 16#08#),
      3546 => to_slv(opcode_type, 16#0C#),
      3547 => to_slv(opcode_type, 16#0F#),
      3548 => to_slv(opcode_type, 16#07#),
      3549 => to_slv(opcode_type, 16#11#),
      3550 => to_slv(opcode_type, 16#0A#),
      3551 to 3551 => (others => '0'),

      -- Program 111...
      3552 => to_slv(opcode_type, 16#07#),
      3553 => to_slv(opcode_type, 16#08#),
      3554 => to_slv(opcode_type, 16#06#),
      3555 => to_slv(opcode_type, 16#07#),
      3556 => to_slv(opcode_type, 16#0E#),
      3557 => to_slv(opcode_type, 16#10#),
      3558 => to_slv(opcode_type, 16#06#),
      3559 => to_slv(opcode_type, 16#0D#),
      3560 => to_slv(opcode_type, 16#0F#),
      3561 => to_slv(opcode_type, 16#07#),
      3562 => to_slv(opcode_type, 16#07#),
      3563 => to_slv(opcode_type, 16#0E#),
      3564 => to_slv(opcode_type, 16#95#),
      3565 => to_slv(opcode_type, 16#09#),
      3566 => to_slv(opcode_type, 16#0B#),
      3567 => to_slv(opcode_type, 16#0C#),
      3568 => to_slv(opcode_type, 16#06#),
      3569 => to_slv(opcode_type, 16#09#),
      3570 => to_slv(opcode_type, 16#08#),
      3571 => to_slv(opcode_type, 16#0A#),
      3572 => to_slv(opcode_type, 16#0E#),
      3573 => to_slv(opcode_type, 16#08#),
      3574 => to_slv(opcode_type, 16#0C#),
      3575 => to_slv(opcode_type, 16#0E#),
      3576 => to_slv(opcode_type, 16#09#),
      3577 => to_slv(opcode_type, 16#09#),
      3578 => to_slv(opcode_type, 16#11#),
      3579 => to_slv(opcode_type, 16#C5#),
      3580 => to_slv(opcode_type, 16#09#),
      3581 => to_slv(opcode_type, 16#0C#),
      3582 => to_slv(opcode_type, 16#64#),
      3583 to 3583 => (others => '0'),

      -- Program 112...
      3584 => to_slv(opcode_type, 16#06#),
      3585 => to_slv(opcode_type, 16#08#),
      3586 => to_slv(opcode_type, 16#09#),
      3587 => to_slv(opcode_type, 16#09#),
      3588 => to_slv(opcode_type, 16#BB#),
      3589 => to_slv(opcode_type, 16#11#),
      3590 => to_slv(opcode_type, 16#06#),
      3591 => to_slv(opcode_type, 16#0C#),
      3592 => to_slv(opcode_type, 16#0A#),
      3593 => to_slv(opcode_type, 16#09#),
      3594 => to_slv(opcode_type, 16#06#),
      3595 => to_slv(opcode_type, 16#11#),
      3596 => to_slv(opcode_type, 16#0A#),
      3597 => to_slv(opcode_type, 16#07#),
      3598 => to_slv(opcode_type, 16#0C#),
      3599 => to_slv(opcode_type, 16#11#),
      3600 => to_slv(opcode_type, 16#07#),
      3601 => to_slv(opcode_type, 16#07#),
      3602 => to_slv(opcode_type, 16#07#),
      3603 => to_slv(opcode_type, 16#B2#),
      3604 => to_slv(opcode_type, 16#AE#),
      3605 => to_slv(opcode_type, 16#09#),
      3606 => to_slv(opcode_type, 16#0A#),
      3607 => to_slv(opcode_type, 16#11#),
      3608 => to_slv(opcode_type, 16#09#),
      3609 => to_slv(opcode_type, 16#06#),
      3610 => to_slv(opcode_type, 16#0A#),
      3611 => to_slv(opcode_type, 16#0D#),
      3612 => to_slv(opcode_type, 16#09#),
      3613 => to_slv(opcode_type, 16#0B#),
      3614 => to_slv(opcode_type, 16#0E#),
      3615 to 3615 => (others => '0'),

      -- Program 113...
      3616 => to_slv(opcode_type, 16#06#),
      3617 => to_slv(opcode_type, 16#08#),
      3618 => to_slv(opcode_type, 16#08#),
      3619 => to_slv(opcode_type, 16#07#),
      3620 => to_slv(opcode_type, 16#0F#),
      3621 => to_slv(opcode_type, 16#0F#),
      3622 => to_slv(opcode_type, 16#06#),
      3623 => to_slv(opcode_type, 16#11#),
      3624 => to_slv(opcode_type, 16#11#),
      3625 => to_slv(opcode_type, 16#08#),
      3626 => to_slv(opcode_type, 16#09#),
      3627 => to_slv(opcode_type, 16#1D#),
      3628 => to_slv(opcode_type, 16#0F#),
      3629 => to_slv(opcode_type, 16#06#),
      3630 => to_slv(opcode_type, 16#0D#),
      3631 => to_slv(opcode_type, 16#0F#),
      3632 => to_slv(opcode_type, 16#09#),
      3633 => to_slv(opcode_type, 16#07#),
      3634 => to_slv(opcode_type, 16#07#),
      3635 => to_slv(opcode_type, 16#0B#),
      3636 => to_slv(opcode_type, 16#10#),
      3637 => to_slv(opcode_type, 16#08#),
      3638 => to_slv(opcode_type, 16#0B#),
      3639 => to_slv(opcode_type, 16#0A#),
      3640 => to_slv(opcode_type, 16#07#),
      3641 => to_slv(opcode_type, 16#08#),
      3642 => to_slv(opcode_type, 16#0D#),
      3643 => to_slv(opcode_type, 16#0D#),
      3644 => to_slv(opcode_type, 16#09#),
      3645 => to_slv(opcode_type, 16#10#),
      3646 => to_slv(opcode_type, 16#0F#),
      3647 to 3647 => (others => '0'),

      -- Program 114...
      3648 => to_slv(opcode_type, 16#08#),
      3649 => to_slv(opcode_type, 16#07#),
      3650 => to_slv(opcode_type, 16#06#),
      3651 => to_slv(opcode_type, 16#09#),
      3652 => to_slv(opcode_type, 16#0D#),
      3653 => to_slv(opcode_type, 16#0B#),
      3654 => to_slv(opcode_type, 16#09#),
      3655 => to_slv(opcode_type, 16#0C#),
      3656 => to_slv(opcode_type, 16#0B#),
      3657 => to_slv(opcode_type, 16#06#),
      3658 => to_slv(opcode_type, 16#07#),
      3659 => to_slv(opcode_type, 16#0E#),
      3660 => to_slv(opcode_type, 16#0D#),
      3661 => to_slv(opcode_type, 16#09#),
      3662 => to_slv(opcode_type, 16#1D#),
      3663 => to_slv(opcode_type, 16#0C#),
      3664 => to_slv(opcode_type, 16#08#),
      3665 => to_slv(opcode_type, 16#07#),
      3666 => to_slv(opcode_type, 16#09#),
      3667 => to_slv(opcode_type, 16#0F#),
      3668 => to_slv(opcode_type, 16#0D#),
      3669 => to_slv(opcode_type, 16#07#),
      3670 => to_slv(opcode_type, 16#0F#),
      3671 => to_slv(opcode_type, 16#0A#),
      3672 => to_slv(opcode_type, 16#08#),
      3673 => to_slv(opcode_type, 16#08#),
      3674 => to_slv(opcode_type, 16#8D#),
      3675 => to_slv(opcode_type, 16#11#),
      3676 => to_slv(opcode_type, 16#06#),
      3677 => to_slv(opcode_type, 16#0B#),
      3678 => to_slv(opcode_type, 16#9E#),
      3679 to 3679 => (others => '0'),

      -- Program 115...
      3680 => to_slv(opcode_type, 16#08#),
      3681 => to_slv(opcode_type, 16#08#),
      3682 => to_slv(opcode_type, 16#07#),
      3683 => to_slv(opcode_type, 16#09#),
      3684 => to_slv(opcode_type, 16#0D#),
      3685 => to_slv(opcode_type, 16#0E#),
      3686 => to_slv(opcode_type, 16#07#),
      3687 => to_slv(opcode_type, 16#0E#),
      3688 => to_slv(opcode_type, 16#0B#),
      3689 => to_slv(opcode_type, 16#08#),
      3690 => to_slv(opcode_type, 16#09#),
      3691 => to_slv(opcode_type, 16#10#),
      3692 => to_slv(opcode_type, 16#11#),
      3693 => to_slv(opcode_type, 16#09#),
      3694 => to_slv(opcode_type, 16#0A#),
      3695 => to_slv(opcode_type, 16#D4#),
      3696 => to_slv(opcode_type, 16#09#),
      3697 => to_slv(opcode_type, 16#08#),
      3698 => to_slv(opcode_type, 16#06#),
      3699 => to_slv(opcode_type, 16#0D#),
      3700 => to_slv(opcode_type, 16#10#),
      3701 => to_slv(opcode_type, 16#06#),
      3702 => to_slv(opcode_type, 16#0A#),
      3703 => to_slv(opcode_type, 16#0A#),
      3704 => to_slv(opcode_type, 16#06#),
      3705 => to_slv(opcode_type, 16#07#),
      3706 => to_slv(opcode_type, 16#11#),
      3707 => to_slv(opcode_type, 16#10#),
      3708 => to_slv(opcode_type, 16#09#),
      3709 => to_slv(opcode_type, 16#11#),
      3710 => to_slv(opcode_type, 16#0F#),
      3711 to 3711 => (others => '0'),

      -- Program 116...
      3712 => to_slv(opcode_type, 16#07#),
      3713 => to_slv(opcode_type, 16#08#),
      3714 => to_slv(opcode_type, 16#07#),
      3715 => to_slv(opcode_type, 16#06#),
      3716 => to_slv(opcode_type, 16#0D#),
      3717 => to_slv(opcode_type, 16#0D#),
      3718 => to_slv(opcode_type, 16#09#),
      3719 => to_slv(opcode_type, 16#0D#),
      3720 => to_slv(opcode_type, 16#9F#),
      3721 => to_slv(opcode_type, 16#07#),
      3722 => to_slv(opcode_type, 16#08#),
      3723 => to_slv(opcode_type, 16#0C#),
      3724 => to_slv(opcode_type, 16#0D#),
      3725 => to_slv(opcode_type, 16#06#),
      3726 => to_slv(opcode_type, 16#0E#),
      3727 => to_slv(opcode_type, 16#0C#),
      3728 => to_slv(opcode_type, 16#06#),
      3729 => to_slv(opcode_type, 16#08#),
      3730 => to_slv(opcode_type, 16#08#),
      3731 => to_slv(opcode_type, 16#0F#),
      3732 => to_slv(opcode_type, 16#0D#),
      3733 => to_slv(opcode_type, 16#07#),
      3734 => to_slv(opcode_type, 16#0B#),
      3735 => to_slv(opcode_type, 16#0B#),
      3736 => to_slv(opcode_type, 16#06#),
      3737 => to_slv(opcode_type, 16#09#),
      3738 => to_slv(opcode_type, 16#1E#),
      3739 => to_slv(opcode_type, 16#0A#),
      3740 => to_slv(opcode_type, 16#08#),
      3741 => to_slv(opcode_type, 16#10#),
      3742 => to_slv(opcode_type, 16#0F#),
      3743 to 3743 => (others => '0'),

      -- Program 117...
      3744 => to_slv(opcode_type, 16#09#),
      3745 => to_slv(opcode_type, 16#06#),
      3746 => to_slv(opcode_type, 16#06#),
      3747 => to_slv(opcode_type, 16#06#),
      3748 => to_slv(opcode_type, 16#0B#),
      3749 => to_slv(opcode_type, 16#0C#),
      3750 => to_slv(opcode_type, 16#07#),
      3751 => to_slv(opcode_type, 16#10#),
      3752 => to_slv(opcode_type, 16#0A#),
      3753 => to_slv(opcode_type, 16#09#),
      3754 => to_slv(opcode_type, 16#06#),
      3755 => to_slv(opcode_type, 16#10#),
      3756 => to_slv(opcode_type, 16#0F#),
      3757 => to_slv(opcode_type, 16#09#),
      3758 => to_slv(opcode_type, 16#10#),
      3759 => to_slv(opcode_type, 16#E8#),
      3760 => to_slv(opcode_type, 16#08#),
      3761 => to_slv(opcode_type, 16#07#),
      3762 => to_slv(opcode_type, 16#07#),
      3763 => to_slv(opcode_type, 16#B2#),
      3764 => to_slv(opcode_type, 16#0B#),
      3765 => to_slv(opcode_type, 16#09#),
      3766 => to_slv(opcode_type, 16#10#),
      3767 => to_slv(opcode_type, 16#0E#),
      3768 => to_slv(opcode_type, 16#06#),
      3769 => to_slv(opcode_type, 16#09#),
      3770 => to_slv(opcode_type, 16#0F#),
      3771 => to_slv(opcode_type, 16#0B#),
      3772 => to_slv(opcode_type, 16#07#),
      3773 => to_slv(opcode_type, 16#0C#),
      3774 => to_slv(opcode_type, 16#0D#),
      3775 to 3775 => (others => '0'),

      -- Program 118...
      3776 => to_slv(opcode_type, 16#09#),
      3777 => to_slv(opcode_type, 16#06#),
      3778 => to_slv(opcode_type, 16#07#),
      3779 => to_slv(opcode_type, 16#07#),
      3780 => to_slv(opcode_type, 16#0C#),
      3781 => to_slv(opcode_type, 16#0F#),
      3782 => to_slv(opcode_type, 16#09#),
      3783 => to_slv(opcode_type, 16#0C#),
      3784 => to_slv(opcode_type, 16#0B#),
      3785 => to_slv(opcode_type, 16#09#),
      3786 => to_slv(opcode_type, 16#06#),
      3787 => to_slv(opcode_type, 16#0A#),
      3788 => to_slv(opcode_type, 16#0C#),
      3789 => to_slv(opcode_type, 16#09#),
      3790 => to_slv(opcode_type, 16#0A#),
      3791 => to_slv(opcode_type, 16#0B#),
      3792 => to_slv(opcode_type, 16#07#),
      3793 => to_slv(opcode_type, 16#07#),
      3794 => to_slv(opcode_type, 16#07#),
      3795 => to_slv(opcode_type, 16#0F#),
      3796 => to_slv(opcode_type, 16#0F#),
      3797 => to_slv(opcode_type, 16#08#),
      3798 => to_slv(opcode_type, 16#0A#),
      3799 => to_slv(opcode_type, 16#0A#),
      3800 => to_slv(opcode_type, 16#08#),
      3801 => to_slv(opcode_type, 16#06#),
      3802 => to_slv(opcode_type, 16#0E#),
      3803 => to_slv(opcode_type, 16#0D#),
      3804 => to_slv(opcode_type, 16#09#),
      3805 => to_slv(opcode_type, 16#0B#),
      3806 => to_slv(opcode_type, 16#10#),
      3807 to 3807 => (others => '0'),

      -- Program 119...
      3808 => to_slv(opcode_type, 16#06#),
      3809 => to_slv(opcode_type, 16#09#),
      3810 => to_slv(opcode_type, 16#09#),
      3811 => to_slv(opcode_type, 16#06#),
      3812 => to_slv(opcode_type, 16#0C#),
      3813 => to_slv(opcode_type, 16#0D#),
      3814 => to_slv(opcode_type, 16#06#),
      3815 => to_slv(opcode_type, 16#11#),
      3816 => to_slv(opcode_type, 16#0C#),
      3817 => to_slv(opcode_type, 16#08#),
      3818 => to_slv(opcode_type, 16#08#),
      3819 => to_slv(opcode_type, 16#0B#),
      3820 => to_slv(opcode_type, 16#0E#),
      3821 => to_slv(opcode_type, 16#06#),
      3822 => to_slv(opcode_type, 16#0A#),
      3823 => to_slv(opcode_type, 16#0C#),
      3824 => to_slv(opcode_type, 16#06#),
      3825 => to_slv(opcode_type, 16#09#),
      3826 => to_slv(opcode_type, 16#09#),
      3827 => to_slv(opcode_type, 16#0A#),
      3828 => to_slv(opcode_type, 16#11#),
      3829 => to_slv(opcode_type, 16#08#),
      3830 => to_slv(opcode_type, 16#0B#),
      3831 => to_slv(opcode_type, 16#0F#),
      3832 => to_slv(opcode_type, 16#06#),
      3833 => to_slv(opcode_type, 16#07#),
      3834 => to_slv(opcode_type, 16#11#),
      3835 => to_slv(opcode_type, 16#0D#),
      3836 => to_slv(opcode_type, 16#08#),
      3837 => to_slv(opcode_type, 16#0B#),
      3838 => to_slv(opcode_type, 16#0C#),
      3839 to 3839 => (others => '0'),

      -- Program 120...
      3840 => to_slv(opcode_type, 16#07#),
      3841 => to_slv(opcode_type, 16#06#),
      3842 => to_slv(opcode_type, 16#08#),
      3843 => to_slv(opcode_type, 16#06#),
      3844 => to_slv(opcode_type, 16#0A#),
      3845 => to_slv(opcode_type, 16#0B#),
      3846 => to_slv(opcode_type, 16#09#),
      3847 => to_slv(opcode_type, 16#0D#),
      3848 => to_slv(opcode_type, 16#0D#),
      3849 => to_slv(opcode_type, 16#08#),
      3850 => to_slv(opcode_type, 16#07#),
      3851 => to_slv(opcode_type, 16#0A#),
      3852 => to_slv(opcode_type, 16#11#),
      3853 => to_slv(opcode_type, 16#06#),
      3854 => to_slv(opcode_type, 16#10#),
      3855 => to_slv(opcode_type, 16#10#),
      3856 => to_slv(opcode_type, 16#09#),
      3857 => to_slv(opcode_type, 16#07#),
      3858 => to_slv(opcode_type, 16#06#),
      3859 => to_slv(opcode_type, 16#11#),
      3860 => to_slv(opcode_type, 16#0B#),
      3861 => to_slv(opcode_type, 16#06#),
      3862 => to_slv(opcode_type, 16#0C#),
      3863 => to_slv(opcode_type, 16#DB#),
      3864 => to_slv(opcode_type, 16#07#),
      3865 => to_slv(opcode_type, 16#08#),
      3866 => to_slv(opcode_type, 16#0B#),
      3867 => to_slv(opcode_type, 16#0C#),
      3868 => to_slv(opcode_type, 16#06#),
      3869 => to_slv(opcode_type, 16#0F#),
      3870 => to_slv(opcode_type, 16#0B#),
      3871 to 3871 => (others => '0'),

      -- Program 121...
      3872 => to_slv(opcode_type, 16#09#),
      3873 => to_slv(opcode_type, 16#09#),
      3874 => to_slv(opcode_type, 16#06#),
      3875 => to_slv(opcode_type, 16#06#),
      3876 => to_slv(opcode_type, 16#0B#),
      3877 => to_slv(opcode_type, 16#10#),
      3878 => to_slv(opcode_type, 16#08#),
      3879 => to_slv(opcode_type, 16#11#),
      3880 => to_slv(opcode_type, 16#0A#),
      3881 => to_slv(opcode_type, 16#08#),
      3882 => to_slv(opcode_type, 16#07#),
      3883 => to_slv(opcode_type, 16#0B#),
      3884 => to_slv(opcode_type, 16#11#),
      3885 => to_slv(opcode_type, 16#08#),
      3886 => to_slv(opcode_type, 16#82#),
      3887 => to_slv(opcode_type, 16#11#),
      3888 => to_slv(opcode_type, 16#07#),
      3889 => to_slv(opcode_type, 16#08#),
      3890 => to_slv(opcode_type, 16#06#),
      3891 => to_slv(opcode_type, 16#22#),
      3892 => to_slv(opcode_type, 16#0E#),
      3893 => to_slv(opcode_type, 16#06#),
      3894 => to_slv(opcode_type, 16#11#),
      3895 => to_slv(opcode_type, 16#0D#),
      3896 => to_slv(opcode_type, 16#07#),
      3897 => to_slv(opcode_type, 16#07#),
      3898 => to_slv(opcode_type, 16#F5#),
      3899 => to_slv(opcode_type, 16#0D#),
      3900 => to_slv(opcode_type, 16#07#),
      3901 => to_slv(opcode_type, 16#0D#),
      3902 => to_slv(opcode_type, 16#0D#),
      3903 to 3903 => (others => '0'),

      -- Program 122...
      3904 => to_slv(opcode_type, 16#09#),
      3905 => to_slv(opcode_type, 16#06#),
      3906 => to_slv(opcode_type, 16#06#),
      3907 => to_slv(opcode_type, 16#09#),
      3908 => to_slv(opcode_type, 16#6F#),
      3909 => to_slv(opcode_type, 16#11#),
      3910 => to_slv(opcode_type, 16#09#),
      3911 => to_slv(opcode_type, 16#11#),
      3912 => to_slv(opcode_type, 16#10#),
      3913 => to_slv(opcode_type, 16#09#),
      3914 => to_slv(opcode_type, 16#07#),
      3915 => to_slv(opcode_type, 16#10#),
      3916 => to_slv(opcode_type, 16#0D#),
      3917 => to_slv(opcode_type, 16#06#),
      3918 => to_slv(opcode_type, 16#0B#),
      3919 => to_slv(opcode_type, 16#0E#),
      3920 => to_slv(opcode_type, 16#07#),
      3921 => to_slv(opcode_type, 16#06#),
      3922 => to_slv(opcode_type, 16#07#),
      3923 => to_slv(opcode_type, 16#0F#),
      3924 => to_slv(opcode_type, 16#11#),
      3925 => to_slv(opcode_type, 16#08#),
      3926 => to_slv(opcode_type, 16#10#),
      3927 => to_slv(opcode_type, 16#0C#),
      3928 => to_slv(opcode_type, 16#06#),
      3929 => to_slv(opcode_type, 16#09#),
      3930 => to_slv(opcode_type, 16#0A#),
      3931 => to_slv(opcode_type, 16#E8#),
      3932 => to_slv(opcode_type, 16#08#),
      3933 => to_slv(opcode_type, 16#60#),
      3934 => to_slv(opcode_type, 16#0C#),
      3935 to 3935 => (others => '0'),

      -- Program 123...
      3936 => to_slv(opcode_type, 16#09#),
      3937 => to_slv(opcode_type, 16#09#),
      3938 => to_slv(opcode_type, 16#06#),
      3939 => to_slv(opcode_type, 16#07#),
      3940 => to_slv(opcode_type, 16#0E#),
      3941 => to_slv(opcode_type, 16#0F#),
      3942 => to_slv(opcode_type, 16#06#),
      3943 => to_slv(opcode_type, 16#0B#),
      3944 => to_slv(opcode_type, 16#0B#),
      3945 => to_slv(opcode_type, 16#06#),
      3946 => to_slv(opcode_type, 16#08#),
      3947 => to_slv(opcode_type, 16#11#),
      3948 => to_slv(opcode_type, 16#0A#),
      3949 => to_slv(opcode_type, 16#07#),
      3950 => to_slv(opcode_type, 16#0C#),
      3951 => to_slv(opcode_type, 16#28#),
      3952 => to_slv(opcode_type, 16#08#),
      3953 => to_slv(opcode_type, 16#09#),
      3954 => to_slv(opcode_type, 16#07#),
      3955 => to_slv(opcode_type, 16#EE#),
      3956 => to_slv(opcode_type, 16#0B#),
      3957 => to_slv(opcode_type, 16#07#),
      3958 => to_slv(opcode_type, 16#0B#),
      3959 => to_slv(opcode_type, 16#0C#),
      3960 => to_slv(opcode_type, 16#09#),
      3961 => to_slv(opcode_type, 16#08#),
      3962 => to_slv(opcode_type, 16#0A#),
      3963 => to_slv(opcode_type, 16#0A#),
      3964 => to_slv(opcode_type, 16#08#),
      3965 => to_slv(opcode_type, 16#10#),
      3966 => to_slv(opcode_type, 16#0F#),
      3967 to 3967 => (others => '0'),

      -- Program 124...
      3968 => to_slv(opcode_type, 16#06#),
      3969 => to_slv(opcode_type, 16#06#),
      3970 => to_slv(opcode_type, 16#06#),
      3971 => to_slv(opcode_type, 16#07#),
      3972 => to_slv(opcode_type, 16#10#),
      3973 => to_slv(opcode_type, 16#0E#),
      3974 => to_slv(opcode_type, 16#07#),
      3975 => to_slv(opcode_type, 16#0A#),
      3976 => to_slv(opcode_type, 16#10#),
      3977 => to_slv(opcode_type, 16#09#),
      3978 => to_slv(opcode_type, 16#09#),
      3979 => to_slv(opcode_type, 16#0B#),
      3980 => to_slv(opcode_type, 16#A4#),
      3981 => to_slv(opcode_type, 16#06#),
      3982 => to_slv(opcode_type, 16#2A#),
      3983 => to_slv(opcode_type, 16#0F#),
      3984 => to_slv(opcode_type, 16#08#),
      3985 => to_slv(opcode_type, 16#08#),
      3986 => to_slv(opcode_type, 16#06#),
      3987 => to_slv(opcode_type, 16#11#),
      3988 => to_slv(opcode_type, 16#0C#),
      3989 => to_slv(opcode_type, 16#09#),
      3990 => to_slv(opcode_type, 16#0D#),
      3991 => to_slv(opcode_type, 16#0C#),
      3992 => to_slv(opcode_type, 16#07#),
      3993 => to_slv(opcode_type, 16#07#),
      3994 => to_slv(opcode_type, 16#E0#),
      3995 => to_slv(opcode_type, 16#0E#),
      3996 => to_slv(opcode_type, 16#06#),
      3997 => to_slv(opcode_type, 16#10#),
      3998 => to_slv(opcode_type, 16#0D#),
      3999 to 3999 => (others => '0'),

      -- Program 125...
      4000 => to_slv(opcode_type, 16#07#),
      4001 => to_slv(opcode_type, 16#07#),
      4002 => to_slv(opcode_type, 16#07#),
      4003 => to_slv(opcode_type, 16#07#),
      4004 => to_slv(opcode_type, 16#0A#),
      4005 => to_slv(opcode_type, 16#0C#),
      4006 => to_slv(opcode_type, 16#08#),
      4007 => to_slv(opcode_type, 16#0F#),
      4008 => to_slv(opcode_type, 16#9C#),
      4009 => to_slv(opcode_type, 16#09#),
      4010 => to_slv(opcode_type, 16#09#),
      4011 => to_slv(opcode_type, 16#0C#),
      4012 => to_slv(opcode_type, 16#0B#),
      4013 => to_slv(opcode_type, 16#09#),
      4014 => to_slv(opcode_type, 16#0A#),
      4015 => to_slv(opcode_type, 16#11#),
      4016 => to_slv(opcode_type, 16#07#),
      4017 => to_slv(opcode_type, 16#08#),
      4018 => to_slv(opcode_type, 16#06#),
      4019 => to_slv(opcode_type, 16#11#),
      4020 => to_slv(opcode_type, 16#10#),
      4021 => to_slv(opcode_type, 16#09#),
      4022 => to_slv(opcode_type, 16#0D#),
      4023 => to_slv(opcode_type, 16#0F#),
      4024 => to_slv(opcode_type, 16#06#),
      4025 => to_slv(opcode_type, 16#08#),
      4026 => to_slv(opcode_type, 16#0C#),
      4027 => to_slv(opcode_type, 16#11#),
      4028 => to_slv(opcode_type, 16#07#),
      4029 => to_slv(opcode_type, 16#11#),
      4030 => to_slv(opcode_type, 16#0F#),
      4031 to 4031 => (others => '0'),

      -- Program 126...
      4032 => to_slv(opcode_type, 16#08#),
      4033 => to_slv(opcode_type, 16#06#),
      4034 => to_slv(opcode_type, 16#07#),
      4035 => to_slv(opcode_type, 16#08#),
      4036 => to_slv(opcode_type, 16#0C#),
      4037 => to_slv(opcode_type, 16#0E#),
      4038 => to_slv(opcode_type, 16#06#),
      4039 => to_slv(opcode_type, 16#10#),
      4040 => to_slv(opcode_type, 16#0D#),
      4041 => to_slv(opcode_type, 16#09#),
      4042 => to_slv(opcode_type, 16#07#),
      4043 => to_slv(opcode_type, 16#0D#),
      4044 => to_slv(opcode_type, 16#0E#),
      4045 => to_slv(opcode_type, 16#08#),
      4046 => to_slv(opcode_type, 16#D8#),
      4047 => to_slv(opcode_type, 16#0C#),
      4048 => to_slv(opcode_type, 16#06#),
      4049 => to_slv(opcode_type, 16#06#),
      4050 => to_slv(opcode_type, 16#06#),
      4051 => to_slv(opcode_type, 16#64#),
      4052 => to_slv(opcode_type, 16#0E#),
      4053 => to_slv(opcode_type, 16#07#),
      4054 => to_slv(opcode_type, 16#10#),
      4055 => to_slv(opcode_type, 16#0F#),
      4056 => to_slv(opcode_type, 16#06#),
      4057 => to_slv(opcode_type, 16#08#),
      4058 => to_slv(opcode_type, 16#0D#),
      4059 => to_slv(opcode_type, 16#0C#),
      4060 => to_slv(opcode_type, 16#07#),
      4061 => to_slv(opcode_type, 16#0D#),
      4062 => to_slv(opcode_type, 16#11#),
      4063 to 4063 => (others => '0'),

      -- Program 127...
      4064 => to_slv(opcode_type, 16#09#),
      4065 => to_slv(opcode_type, 16#07#),
      4066 => to_slv(opcode_type, 16#06#),
      4067 => to_slv(opcode_type, 16#09#),
      4068 => to_slv(opcode_type, 16#0E#),
      4069 => to_slv(opcode_type, 16#57#),
      4070 => to_slv(opcode_type, 16#09#),
      4071 => to_slv(opcode_type, 16#0F#),
      4072 => to_slv(opcode_type, 16#0B#),
      4073 => to_slv(opcode_type, 16#09#),
      4074 => to_slv(opcode_type, 16#08#),
      4075 => to_slv(opcode_type, 16#11#),
      4076 => to_slv(opcode_type, 16#10#),
      4077 => to_slv(opcode_type, 16#07#),
      4078 => to_slv(opcode_type, 16#11#),
      4079 => to_slv(opcode_type, 16#0F#),
      4080 => to_slv(opcode_type, 16#09#),
      4081 => to_slv(opcode_type, 16#08#),
      4082 => to_slv(opcode_type, 16#09#),
      4083 => to_slv(opcode_type, 16#0D#),
      4084 => to_slv(opcode_type, 16#6F#),
      4085 => to_slv(opcode_type, 16#06#),
      4086 => to_slv(opcode_type, 16#11#),
      4087 => to_slv(opcode_type, 16#0C#),
      4088 => to_slv(opcode_type, 16#06#),
      4089 => to_slv(opcode_type, 16#08#),
      4090 => to_slv(opcode_type, 16#10#),
      4091 => to_slv(opcode_type, 16#10#),
      4092 => to_slv(opcode_type, 16#08#),
      4093 => to_slv(opcode_type, 16#E3#),
      4094 => to_slv(opcode_type, 16#0B#),
      4095 to 4095 => (others => '0')
  )
);

end package;